library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;
use ieee.numeric_std.all;

entity spaceship is
    Port (
        address : in STD_LOGIC_VECTOR(14 downto 0);
        data_out : out STD_LOGIC_VECTOR(23 downto 0)
    );
end entity spaceship;

architecture Behavioral of spaceship is
    type ROM_Type is array (0 to 22499) of STD_LOGIC_VECTOR(23 downto 0);
    constant ROM_Data : ROM_Type := (
0 => "000000000000000000000000",
1 => "000000000000000000000000",
2 => "000000000000000000000000",
3 => "000000000000000000000000",
4 => "000000000000000000000000",
5 => "000000000000000000000000",
6 => "000000000000000000000000",
7 => "000000000000000000000000",
8 => "000000000000000000000000",
9 => "000000000000000000000000",
10 => "000000000000000000000000",
11 => "000000000000000000000000",
12 => "000000000000000000000000",
13 => "000000000000000000000000",
14 => "000000000000000000000000",
15 => "000000000000000000000000",
16 => "000000000000000000000000",
17 => "000000000000000000000000",
18 => "000000000000000000000000",
19 => "000000000000000000000000",
20 => "000000000000000000000000",
21 => "000000000000000000000000",
22 => "000000000000000000000000",
23 => "000000000000000000000000",
24 => "000000000000000000000000",
25 => "000000000000000000000000",
26 => "000000000000000000000000",
27 => "000000000000000000000000",
28 => "000000000000000000000000",
29 => "000000000000000000000000",
30 => "000000000000000000000000",
31 => "000000000000000000000000",
32 => "000000000000000000000000",
33 => "000000000000000000000000",
34 => "000000000000000000000000",
35 => "000000000000000000000000",
36 => "000000000000000000000000",
37 => "000000000000000000000000",
38 => "000000000000000000000000",
39 => "000000000000000000000000",
40 => "000000000000000000000000",
41 => "000000000000000000000000",
42 => "000000000000000000000000",
43 => "000000000000000000000000",
44 => "000000000000000000000000",
45 => "000000000000000000000000",
46 => "000000000000000000000000",
47 => "000000000000000000000000",
48 => "000000000000000000000000",
49 => "000000000000000000000000",
50 => "000000000000000000000000",
51 => "000000000000000000000000",
52 => "000000000000000000000000",
53 => "000000000000000000000000",
54 => "000000000000000000000000",
55 => "000000000000000000000000",
56 => "000000000000000000000000",
57 => "000000000000000000000000",
58 => "000000000000000000000000",
59 => "000000000000000000000000",
60 => "000000000000000000000000",
61 => "000000000000000000000000",
62 => "000000000000000000000000",
63 => "000000000000000000000000",
64 => "000000000000000000000000",
65 => "000000000000000000000000",
66 => "000000000000000000000000",
67 => "000000000000000000000000",
68 => "000000000000000000000000",
69 => "000000000000000000000000",
70 => "000000000000000000000000",
71 => "000000000000000000000000",
72 => "000000000000000000000000",
73 => "000000000000000000000000",
74 => "000000000000000000000000",
75 => "000000000000000000000000",
76 => "000000000000000000000000",
77 => "000000000000000000000000",
78 => "000000000000000000000000",
79 => "000000000000000000000000",
80 => "000000000000000000000000",
81 => "000000000000000000000000",
82 => "000000000000000000000000",
83 => "000000000000000000000000",
84 => "000000000000000000000000",
85 => "000000000000000000000000",
86 => "000000000000000000000000",
87 => "000000000000000000000000",
88 => "000000000000000000000000",
89 => "000000000000000000000000",
90 => "000000000000000000000000",
91 => "000000000000000000000000",
92 => "000000000000000000000000",
93 => "000000000000000000000000",
94 => "000000000000000000000000",
95 => "000000000000000000000000",
96 => "000000000000000000000000",
97 => "000000000000000000000000",
98 => "000000000000000000000000",
99 => "000000000000000000000000",
100 => "000000000000000000000000",
101 => "000000000000000000000000",
102 => "000000000000000000000000",
103 => "000000000000000000000000",
104 => "000000000000000000000000",
105 => "000000000000000000000000",
106 => "000000000000000000000000",
107 => "000000000000000000000000",
108 => "000000000000000000000000",
109 => "000000000000000000000000",
110 => "000000000000000000000000",
111 => "000000000000000000000000",
112 => "000000000000000000000000",
113 => "000000000000000000000000",
114 => "000000000000000000000000",
115 => "000000000000000000000000",
116 => "000000000000000000000000",
117 => "000000000000000000000000",
118 => "000000000000000000000000",
119 => "000000000000000000000000",
120 => "000000000000000000000000",
121 => "000000000000000000000000",
122 => "000000000000000000000000",
123 => "000000000000000000000000",
124 => "000000000000000000000000",
125 => "000000000000000000000000",
126 => "000000000000000000000000",
127 => "000000000000000000000000",
128 => "000000000000000000000000",
129 => "000000000000000000000000",
130 => "000000000000000000000000",
131 => "000000000000000000000000",
132 => "000000000000000000000000",
133 => "000000000000000000000000",
134 => "000000000000000000000000",
135 => "000000000000000000000000",
136 => "000000000000000000000000",
137 => "000000000000000000000000",
138 => "000000000000000000000000",
139 => "000000000000000000000000",
140 => "000000000000000000000000",
141 => "000000000000000000000000",
142 => "000000000000000000000000",
143 => "000000000000000000000000",
144 => "000000000000000000000000",
145 => "000000000000000000000000",
146 => "000000000000000000000000",
147 => "000000000000000000000000",
148 => "000000000000000000000000",
149 => "000000000000000000000000",
150 => "000000000000000000000000",
151 => "000000000000000000000000",
152 => "000000000000000000000000",
153 => "000000000000000000000000",
154 => "000000000000000000000000",
155 => "000000000000000000000000",
156 => "000000000000000000000000",
157 => "000000000000000000000000",
158 => "000000000000000000000000",
159 => "000000000000000000000000",
160 => "000000000000000000000000",
161 => "000000000000000000000000",
162 => "000000000000000000000000",
163 => "000000000000000000000000",
164 => "000000000000000000000000",
165 => "000000000000000000000000",
166 => "000000000000000000000000",
167 => "000000000000000000000000",
168 => "000000000000000000000000",
169 => "000000000000000000000000",
170 => "000000000000000000000000",
171 => "000000000000000000000000",
172 => "000000000000000000000000",
173 => "000000000000000000000000",
174 => "000000000000000000000000",
175 => "000000000000000000000000",
176 => "000000000000000000000000",
177 => "000000000000000000000000",
178 => "000000000000000000000000",
179 => "000000000000000000000000",
180 => "000000000000000000000000",
181 => "000000000000000000000000",
182 => "000000000000000000000000",
183 => "000000000000000000000000",
184 => "000000000000000000000000",
185 => "000000000000000000000000",
186 => "000000000000000000000000",
187 => "000000000000000000000000",
188 => "000000000000000000000000",
189 => "000000000000000000000000",
190 => "000000000000000000000000",
191 => "000000000000000000000000",
192 => "000000000000000000000000",
193 => "000000000000000000000000",
194 => "000000000000000000000000",
195 => "000000000000000000000000",
196 => "000000000000000000000000",
197 => "000000000000000000000000",
198 => "000000000000000000000000",
199 => "000000000000000000000000",
200 => "000000000000000000000000",
201 => "000000000000000000000000",
202 => "000000000000000000000000",
203 => "000000000000000000000000",
204 => "000000000000000000000000",
205 => "000000000000000000000000",
206 => "000000000000000000000000",
207 => "000000000000000000000000",
208 => "000000000000000000000000",
209 => "000000000000000000000000",
210 => "000000000000000000000000",
211 => "000000000000000000000000",
212 => "000000000000000000000000",
213 => "000000000000000000000000",
214 => "000000000000000000000000",
215 => "000000000000000000000000",
216 => "000000000000000000000000",
217 => "000000000000000000000000",
218 => "000000000000000000000000",
219 => "000000000000000000000000",
220 => "000000000000000000000000",
221 => "000000000000000000000000",
222 => "000000000000000000000000",
223 => "000000000000000000000000",
224 => "000000000000000000000000",
225 => "000000000000000000000000",
226 => "000000000000000000000000",
227 => "000000000000000000000000",
228 => "000000000000000000000000",
229 => "000000000000000000000000",
230 => "000000000000000000000000",
231 => "000000000000000000000000",
232 => "000000000000000000000000",
233 => "000000000000000000000000",
234 => "000000000000000000000000",
235 => "000000000000000000000000",
236 => "000000000000000000000000",
237 => "000000000000000000000000",
238 => "000000000000000000000000",
239 => "000000000000000000000000",
240 => "000000000000000000000000",
241 => "000000000000000000000000",
242 => "000000000000000000000000",
243 => "000000000000000000000000",
244 => "000000000000000000000000",
245 => "000000000000000000000000",
246 => "000000000000000000000000",
247 => "000000000000000000000000",
248 => "000000000000000000000000",
249 => "000000000000000000000000",
250 => "000000000000000000000000",
251 => "000000000000000000000000",
252 => "000000000000000000000000",
253 => "000000000000000000000000",
254 => "000000000000000000000000",
255 => "000000000000000000000000",
256 => "000000000000000000000000",
257 => "000000000000000000000000",
258 => "000000000000000000000000",
259 => "000000000000000000000000",
260 => "000000000000000000000000",
261 => "000000000000000000000000",
262 => "000000000000000000000000",
263 => "000000000000000000000000",
264 => "000000000000000000000000",
265 => "000000000000000000000000",
266 => "000000000000000000000000",
267 => "000000000000000000000000",
268 => "000000000000000000000000",
269 => "000000000000000000000000",
270 => "000000000000000000000000",
271 => "000000000000000000000000",
272 => "000000000000000000000000",
273 => "000000000000000000000000",
274 => "000000000000000000000000",
275 => "000000000000000000000000",
276 => "000000000000000000000000",
277 => "000000000000000000000000",
278 => "000000000000000000000000",
279 => "000000000000000000000000",
280 => "000000000000000000000000",
281 => "000000000000000000000000",
282 => "000000000000000000000000",
283 => "000000000000000000000000",
284 => "000000000000000000000000",
285 => "000000000000000000000000",
286 => "000000000000000000000000",
287 => "000000000000000000000000",
288 => "000000000000000000000000",
289 => "000000000000000000000000",
290 => "000000000000000000000000",
291 => "000000000000000000000000",
292 => "000000000000000000000000",
293 => "000000000000000000000000",
294 => "000000000000000000000000",
295 => "000000000000000000000000",
296 => "000000000000000000000000",
297 => "000000000000000000000000",
298 => "000000000000000000000000",
299 => "000000000000000000000000",
300 => "000000000000000000000000",
301 => "000000000000000000000000",
302 => "000000000000000000000000",
303 => "000000000000000000000000",
304 => "000000000000000000000000",
305 => "000000000000000000000000",
306 => "000000000000000000000000",
307 => "000000000000000000000000",
308 => "000000000000000000000000",
309 => "000000000000000000000000",
310 => "000000000000000000000000",
311 => "000000000000000000000000",
312 => "000000000000000000000000",
313 => "000000000000000000000000",
314 => "000000000000000000000000",
315 => "000000000000000000000000",
316 => "000000000000000000000000",
317 => "000000000000000000000000",
318 => "000000000000000000000000",
319 => "000000000000000000000000",
320 => "000000000000000000000000",
321 => "000000000000000000000000",
322 => "000000000000000000000000",
323 => "000000000000000000000000",
324 => "000000000000000000000000",
325 => "000000000000000000000000",
326 => "000000000000000000000000",
327 => "000000000000000000000000",
328 => "000000000000000000000000",
329 => "000000000000000000000000",
330 => "000000000000000000000000",
331 => "000000000000000000000000",
332 => "000000000000000000000000",
333 => "000000000000000000000000",
334 => "000000000000000000000000",
335 => "000000000000000000000000",
336 => "000000000000000000000000",
337 => "000000000000000000000000",
338 => "000000000000000000000000",
339 => "000000000000000000000000",
340 => "000000000000000000000000",
341 => "000000000000000000000000",
342 => "000000000000000000000000",
343 => "000000000000000000000000",
344 => "000000000000000000000000",
345 => "000000000000000000000000",
346 => "000000000000000000000000",
347 => "000000000000000000000000",
348 => "000000000000000000000000",
349 => "000000000000000000000000",
350 => "000000000000000000000000",
351 => "000000000000000000000000",
352 => "000000000000000000000000",
353 => "000000000000000000000000",
354 => "000000000000000000000000",
355 => "000000000000000000000000",
356 => "000000000000000000000000",
357 => "000000000000000000000000",
358 => "000000000000000000000000",
359 => "000000000000000000000000",
360 => "000000000000000000000000",
361 => "000000000000000000000000",
362 => "000000000000000000000000",
363 => "000000000000000000000000",
364 => "000000000000000000000000",
365 => "000000000000000000000000",
366 => "000000000000000000000000",
367 => "000000000000000000000000",
368 => "000000000000000000000000",
369 => "000000000000000000000000",
370 => "000000000000000000000000",
371 => "000000000000000000000000",
372 => "000000000000000000000000",
373 => "000000000000000000000000",
374 => "000000000000000000000000",
375 => "000000000000000000000000",
376 => "000000000000000000000000",
377 => "000000000000000000000000",
378 => "000000000000000000000000",
379 => "000000000000000000000000",
380 => "000000000000000000000000",
381 => "000000000000000000000000",
382 => "000000000000000000000000",
383 => "000000000000000000000000",
384 => "000000000000000000000000",
385 => "000000000000000000000000",
386 => "000000000000000000000000",
387 => "000000000000000000000000",
388 => "000000000000000000000000",
389 => "000000000000000000000000",
390 => "000000000000000000000000",
391 => "000000000000000000000000",
392 => "000000000000000000000000",
393 => "000000000000000000000000",
394 => "000000000000000000000000",
395 => "000000000000000000000000",
396 => "000000000000000000000000",
397 => "000000000000000000000000",
398 => "000000000000000000000000",
399 => "000000000000000000000000",
400 => "000000000000000000000000",
401 => "000000000000000000000000",
402 => "000000000000000000000000",
403 => "000000000000000000000000",
404 => "000000000000000000000000",
405 => "000000000000000000000000",
406 => "000000000000000000000000",
407 => "000000000000000000000000",
408 => "000000000000000000000000",
409 => "000000000000000000000000",
410 => "000000000000000000000000",
411 => "000000000000000000000000",
412 => "000000000000000000000000",
413 => "000000000000000000000000",
414 => "000000000000000000000000",
415 => "000000000000000000000000",
416 => "000000000000000000000000",
417 => "000000000000000000000000",
418 => "000000000000000000000000",
419 => "000000000000000000000000",
420 => "000000000000000000000000",
421 => "000000000000000000000000",
422 => "000000000000000000000000",
423 => "000000000000000000000000",
424 => "000000000000000000000000",
425 => "000000000000000000000000",
426 => "000000000000000000000000",
427 => "000000000000000000000000",
428 => "000000000000000000000000",
429 => "000000000000000000000000",
430 => "000000000000000000000000",
431 => "000000000000000000000000",
432 => "000000000000000000000000",
433 => "000000000000000000000000",
434 => "000000000000000000000000",
435 => "000000000000000000000000",
436 => "000000000000000000000000",
437 => "000000000000000000000000",
438 => "000000000000000000000000",
439 => "000000000000000000000000",
440 => "000000000000000000000000",
441 => "000000000000000000000000",
442 => "000000000000000000000000",
443 => "000000000000000000000000",
444 => "000000000000000000000000",
445 => "000000000000000000000000",
446 => "000000000000000000000000",
447 => "000000000000000000000000",
448 => "000000000000000000000000",
449 => "000000000000000000000000",
450 => "000000000000000000000000",
451 => "000000000000000000000000",
452 => "000000000000000000000000",
453 => "000000000000000000000000",
454 => "000000000000000000000000",
455 => "000000000000000000000000",
456 => "000000000000000000000000",
457 => "000000000000000000000000",
458 => "000000000000000000000000",
459 => "000000000000000000000000",
460 => "000000000000000000000000",
461 => "000000000000000000000000",
462 => "000000000000000000000000",
463 => "000000000000000000000000",
464 => "000000000000000000000000",
465 => "000000000000000000000000",
466 => "000000000000000000000000",
467 => "000000000000000000000000",
468 => "000000000000000000000000",
469 => "000000000000000000000000",
470 => "000000000000000000000000",
471 => "000000000000000000000000",
472 => "000000000000000000000000",
473 => "000000000000000000000000",
474 => "000000000000000000000000",
475 => "000000000000000000000000",
476 => "000000000000000000000000",
477 => "000000000000000000000000",
478 => "000000000000000000000000",
479 => "000000000000000000000000",
480 => "000000000000000000000000",
481 => "000000000000000000000000",
482 => "000000000000000000000000",
483 => "000000000000000000000000",
484 => "000000000000000000000000",
485 => "000000000000000000000000",
486 => "000000000000000000000000",
487 => "000000000000000000000000",
488 => "000000000000000000000000",
489 => "000000000000000000000000",
490 => "000000000000000000000000",
491 => "000000000000000000000000",
492 => "000000000000000000000000",
493 => "000000000000000000000000",
494 => "000000000000000000000000",
495 => "000000000000000000000000",
496 => "000000000000000000000000",
497 => "000000000000000000000000",
498 => "000000000000000000000000",
499 => "000000000000000000000000",
500 => "000000000000000000000000",
501 => "000000000000000000000000",
502 => "000000000000000000000000",
503 => "000000000000000000000000",
504 => "000000000000000000000000",
505 => "000000000000000000000000",
506 => "000000000000000000000000",
507 => "000000000000000000000000",
508 => "000000000000000000000000",
509 => "000000000000000000000000",
510 => "000000000000000000000000",
511 => "000000000000000000000000",
512 => "000000000000000000000000",
513 => "000000000000000000000000",
514 => "000000000000000000000000",
515 => "000000000000000000000000",
516 => "000000000000000000000000",
517 => "000000000000000000000000",
518 => "000000000000000000000000",
519 => "000000000000000000000000",
520 => "000000000000000000000000",
521 => "000000000000000000000000",
522 => "000000000000000000000000",
523 => "000000000000000000000000",
524 => "000000000000000000000000",
525 => "000000000000000000000000",
526 => "000000000000000000000000",
527 => "000000000000000000000000",
528 => "000000000000000000000000",
529 => "000000000000000000000000",
530 => "000000000000000000000000",
531 => "000000000000000000000000",
532 => "000000000000000000000000",
533 => "000000000000000000000000",
534 => "000000000000000000000000",
535 => "000000000000000000000000",
536 => "000000000000000000000000",
537 => "000000000000000000000000",
538 => "000000000000000000000000",
539 => "000000000000000000000000",
540 => "000000000000000000000000",
541 => "000000000000000000000000",
542 => "000000000000000000000000",
543 => "000000000000000000000000",
544 => "000000000000000000000000",
545 => "000000000000000000000000",
546 => "000000000000000000000000",
547 => "000000000000000000000000",
548 => "000000000000000000000000",
549 => "000000000000000000000000",
550 => "000000000000000000000000",
551 => "000000000000000000000000",
552 => "000000000000000000000000",
553 => "000000000000000000000000",
554 => "000000000000000000000000",
555 => "000000000000000000000000",
556 => "000000000000000000000000",
557 => "000000000000000000000000",
558 => "000000000000000000000000",
559 => "000000000000000000000000",
560 => "000000000000000000000000",
561 => "000000000000000000000000",
562 => "000000000000000000000000",
563 => "000000000000000000000000",
564 => "000000000000000000000000",
565 => "000000000000000000000000",
566 => "000000000000000000000000",
567 => "000000000000000000000000",
568 => "000000000000000000000000",
569 => "000000000000000000000000",
570 => "000000000000000000000000",
571 => "000000000000000000000000",
572 => "000000000000000000000000",
573 => "000000000000000000000000",
574 => "000000000000000000000000",
575 => "000000000000000000000000",
576 => "000000000000000000000000",
577 => "000000000000000000000000",
578 => "000000000000000000000000",
579 => "000000000000000000000000",
580 => "000000000000000000000000",
581 => "000000000000000000000000",
582 => "000000000000000000000000",
583 => "000000000000000000000000",
584 => "000000000000000000000000",
585 => "000000000000000000000000",
586 => "000000000000000000000000",
587 => "000000000000000000000000",
588 => "000000000000000000000000",
589 => "000000000000000000000000",
590 => "000000000000000000000000",
591 => "000000000000000000000000",
592 => "000000000000000000000000",
593 => "000000000000000000000000",
594 => "000000000000000000000000",
595 => "000000000000000000000000",
596 => "000000000000000000000000",
597 => "000000000000000000000000",
598 => "000000000000000000000000",
599 => "000000000000000000000000",
600 => "000000000000000000000000",
601 => "000000000000000000000000",
602 => "000000000000000000000000",
603 => "000000000000000000000000",
604 => "000000000000000000000000",
605 => "000000000000000000000000",
606 => "000000000000000000000000",
607 => "000000000000000000000000",
608 => "000000000000000000000000",
609 => "000000000000000000000000",
610 => "000000000000000000000000",
611 => "000000000000000000000000",
612 => "000000000000000000000000",
613 => "000000000000000000000000",
614 => "000000000000000000000000",
615 => "000000000000000000000000",
616 => "000000000000000000000000",
617 => "000000000000000000000000",
618 => "000000000000000000000000",
619 => "000000000000000000000000",
620 => "000000000000000000000000",
621 => "000000000000000000000000",
622 => "000000000000000000000000",
623 => "000000000000000000000000",
624 => "000000000000000000000000",
625 => "000000000000000000000000",
626 => "000000000000000000000000",
627 => "000000000000000000000000",
628 => "000000000000000000000000",
629 => "000000000000000000000000",
630 => "000000000000000000000000",
631 => "000000000000000000000000",
632 => "000000000000000000000000",
633 => "000000000000000000000000",
634 => "000000000000000000000000",
635 => "000000000000000000000000",
636 => "000000000000000000000000",
637 => "000000000000000000000000",
638 => "000000000000000000000000",
639 => "000000000000000000000000",
640 => "000000000000000000000000",
641 => "000000000000000000000000",
642 => "000000000000000000000000",
643 => "000000000000000000000000",
644 => "000000000000000000000000",
645 => "000000000000000000000000",
646 => "000000000000000000000000",
647 => "000000000000000000000000",
648 => "000000000000000000000000",
649 => "000000000000000000000000",
650 => "000000000000000000000000",
651 => "000000000000000000000000",
652 => "000000000000000000000000",
653 => "000000000000000000000000",
654 => "000000000000000000000000",
655 => "000000000000000000000000",
656 => "000000000000000000000000",
657 => "000000000000000000000000",
658 => "000000000000000000000000",
659 => "000000000000000000000000",
660 => "000000000000000000000000",
661 => "000000000000000000000000",
662 => "000000000000000000000000",
663 => "000000000000000000000000",
664 => "000000000000000000000000",
665 => "000000000000000000000000",
666 => "000000000000000000000000",
667 => "000000000000000000000000",
668 => "000000000000000000000000",
669 => "000000000000000000000000",
670 => "000000000000000000000000",
671 => "000000000000000000000000",
672 => "000000000000000000000000",
673 => "000000000000000000000000",
674 => "000000000000000000000000",
675 => "000000000000000000000000",
676 => "000000000000000000000000",
677 => "000000000000000000000000",
678 => "000000000000000000000000",
679 => "000000000000000000000000",
680 => "000000000000000000000000",
681 => "000000000000000000000000",
682 => "000000000000000000000000",
683 => "000000000000000000000000",
684 => "000000000000000000000000",
685 => "000000000000000000000000",
686 => "000000000000000000000000",
687 => "000000000000000000000000",
688 => "000000000000000000000000",
689 => "000000000000000000000000",
690 => "000000000000000000000000",
691 => "000000000000000000000000",
692 => "000000000000000000000000",
693 => "000000000000000000000000",
694 => "000000000000000000000000",
695 => "000000000000000000000000",
696 => "000000000000000000000000",
697 => "000000000000000000000000",
698 => "000000000000000000000000",
699 => "000000000000000000000000",
700 => "000000000000000000000000",
701 => "000000000000000000000000",
702 => "000000000000000000000000",
703 => "000000000000000000000000",
704 => "000000000000000000000000",
705 => "000000000000000000000000",
706 => "000000000000000000000000",
707 => "000000000000000000000000",
708 => "000000000000000000000000",
709 => "000000000000000000000000",
710 => "000000000000000000000000",
711 => "000000000000000000000000",
712 => "000000000000000000000000",
713 => "000000000000000000000000",
714 => "000000000000000000000000",
715 => "000000000000000000000000",
716 => "000000000000000000000000",
717 => "000000000000000000000000",
718 => "000000000000000000000000",
719 => "000000000000000000000000",
720 => "000000000000000000000000",
721 => "000000000000000000000000",
722 => "000000000000000000000000",
723 => "000000000000000000000000",
724 => "000000000000000000000000",
725 => "000000000000000000000000",
726 => "000000000000000000000000",
727 => "000000000000000000000000",
728 => "000000000000000000000000",
729 => "000000000000000000000000",
730 => "000000000000000000000000",
731 => "000000000000000000000000",
732 => "000000000000000000000000",
733 => "000000000000000000000000",
734 => "000000000000000000000000",
735 => "000000000000000000000000",
736 => "000000000000000000000000",
737 => "000000000000000000000000",
738 => "000000000000000000000000",
739 => "000000000000000000000000",
740 => "000000000000000000000000",
741 => "000000000000000000000000",
742 => "000000000000000000000000",
743 => "000000000000000000000000",
744 => "000000000000000000000000",
745 => "000000000000000000000000",
746 => "000000000000000000000000",
747 => "000000000000000000000000",
748 => "000000000000000000000000",
749 => "000000000000000000000000",
750 => "000000000000000000000000",
751 => "000000000000000000000000",
752 => "000000000000000000000000",
753 => "000000000000000000000000",
754 => "000000000000000000000000",
755 => "000000000000000000000000",
756 => "000000000000000000000000",
757 => "000000000000000000000000",
758 => "000000000000000000000000",
759 => "000000000000000000000000",
760 => "000000000000000000000000",
761 => "000000000000000000000000",
762 => "000000000000000000000000",
763 => "000000000000000000000000",
764 => "000000000000000000000000",
765 => "000000000000000000000000",
766 => "000000000000000000000000",
767 => "000000000000000000000000",
768 => "000000000000000000000000",
769 => "000000000000000000000000",
770 => "000000000000000000000000",
771 => "000000000000000000000000",
772 => "000000000000000000000000",
773 => "000000000000000000000000",
774 => "000000000000000000000000",
775 => "000000000000000000000000",
776 => "000000000000000000000000",
777 => "000000000000000000000000",
778 => "000000000000000000000000",
779 => "000000000000000000000000",
780 => "000000000000000000000000",
781 => "000000000000000000000000",
782 => "000000000000000000000000",
783 => "000000000000000000000000",
784 => "000000000000000000000000",
785 => "000000000000000000000000",
786 => "000000000000000000000000",
787 => "000000000000000000000000",
788 => "000000000000000000000000",
789 => "000000000000000000000000",
790 => "000000000000000000000000",
791 => "000000000000000000000000",
792 => "000000000000000000000000",
793 => "000000000000000000000000",
794 => "000000000000000000000000",
795 => "000000000000000000000000",
796 => "000000000000000000000000",
797 => "000000000000000000000000",
798 => "000000000000000000000000",
799 => "000000000000000000000000",
800 => "000000000000000000000000",
801 => "000000000000000000000000",
802 => "000000000000000000000000",
803 => "000000000000000000000000",
804 => "000000000000000000000000",
805 => "000000000000000000000000",
806 => "000000000000000000000000",
807 => "000000000000000000000000",
808 => "000000000000000000000000",
809 => "000000000000000000000000",
810 => "000000000000000000000000",
811 => "000000000000000000000000",
812 => "000000000000000000000000",
813 => "000000000000000000000000",
814 => "000000000000000000000000",
815 => "000000000000000000000000",
816 => "000000000000000000000000",
817 => "000000000000000000000000",
818 => "000000000000000000000000",
819 => "000000000000000000000000",
820 => "000000000000000000000000",
821 => "000000000000000000000000",
822 => "000000000000000000000000",
823 => "000000000000000000000000",
824 => "000000000000000000000000",
825 => "000000000000000000000000",
826 => "000000000000000000000000",
827 => "000000000000000000000000",
828 => "000000000000000000000000",
829 => "000000000000000000000000",
830 => "000000000000000000000000",
831 => "000000000000000000000000",
832 => "000000000000000000000000",
833 => "000000000000000000000000",
834 => "000000000000000000000000",
835 => "000000000000000000000000",
836 => "000000000000000000000000",
837 => "000000000000000000000000",
838 => "000000000000000000000000",
839 => "000000000000000000000000",
840 => "000000000000000000000000",
841 => "000000000000000000000000",
842 => "000000000000000000000000",
843 => "000000000000000000000000",
844 => "000000000000000000000000",
845 => "000000000000000000000000",
846 => "000000000000000000000000",
847 => "000000000000000000000000",
848 => "000000000000000000000000",
849 => "000000000000000000000000",
850 => "000000000000000000000000",
851 => "000000000000000000000000",
852 => "000000000000000000000000",
853 => "000000000000000000000000",
854 => "000000000000000000000000",
855 => "000000000000000000000000",
856 => "000000000000000000000000",
857 => "000000000000000000000000",
858 => "000000000000000000000000",
859 => "000000000000000000000000",
860 => "000000000000000000000000",
861 => "000000000000000000000000",
862 => "000000000000000000000000",
863 => "000000000000000000000000",
864 => "000000000000000000000000",
865 => "000000000000000000000000",
866 => "000000000000000000000000",
867 => "000000000000000000000000",
868 => "000000000000000000000000",
869 => "000000000000000000000000",
870 => "000000000000000000000000",
871 => "000000000000000000000000",
872 => "000000000000000000000000",
873 => "000000000000000000000000",
874 => "000000000000000000000000",
875 => "000000000000000000000000",
876 => "000000000000000000000000",
877 => "000000000000000000000000",
878 => "000000000000000000000000",
879 => "000000000000000000000000",
880 => "000000000000000000000000",
881 => "000000000000000000000000",
882 => "000000000000000000000000",
883 => "000000000000000000000000",
884 => "000000000000000000000000",
885 => "000000000000000000000000",
886 => "000000000000000000000000",
887 => "000000000000000000000000",
888 => "000000000000000000000000",
889 => "000000000000000000000000",
890 => "000000000000000000000000",
891 => "000000000000000000000000",
892 => "000000000000000000000000",
893 => "000000000000000000000000",
894 => "000000000000000000000000",
895 => "000000000000000000000000",
896 => "000000000000000000000000",
897 => "000000000000000000000000",
898 => "000000000000000000000000",
899 => "000000000000000000000000",
900 => "000000000000000000000000",
901 => "000000000000000000000000",
902 => "000000000000000000000000",
903 => "000000000000000000000000",
904 => "000000000000000000000000",
905 => "000000000000000000000000",
906 => "000000000000000000000000",
907 => "000000000000000000000000",
908 => "000000000000000000000000",
909 => "000000000000000000000000",
910 => "000000000000000000000000",
911 => "000000000000000000000000",
912 => "000000000000000000000000",
913 => "000000000000000000000000",
914 => "000000000000000000000000",
915 => "000000000000000000000000",
916 => "000000000000000000000000",
917 => "000000000000000000000000",
918 => "000000000000000000000000",
919 => "000000000000000000000000",
920 => "000000000000000000000000",
921 => "000000000000000000000000",
922 => "000000000000000000000000",
923 => "000000000000000000000000",
924 => "000000000000000000000000",
925 => "000000000000000000000000",
926 => "000000000000000000000000",
927 => "000000000000000000000000",
928 => "000000000000000000000000",
929 => "000000000000000000000000",
930 => "000000000000000000000000",
931 => "000000000000000000000000",
932 => "000000000000000000000000",
933 => "000000000000000000000000",
934 => "000000000000000000000000",
935 => "000000000000000000000000",
936 => "000000000000000000000000",
937 => "000000000000000000000000",
938 => "000000000000000000000000",
939 => "000000000000000000000000",
940 => "000000000000000000000000",
941 => "000000000000000000000000",
942 => "000000000000000000000000",
943 => "000000000000000000000000",
944 => "000000000000000000000000",
945 => "000000000000000000000000",
946 => "000000000000000000000000",
947 => "000000000000000000000000",
948 => "000000000000000000000000",
949 => "000000000000000000000000",
950 => "000000000000000000000000",
951 => "000000000000000000000000",
952 => "000000000000000000000000",
953 => "000000000000000000000000",
954 => "000000000000000000000000",
955 => "000000000000000000000000",
956 => "000000000000000000000000",
957 => "000000000000000000000000",
958 => "000000000000000000000000",
959 => "000000000000000000000000",
960 => "000000000000000000000000",
961 => "000000000000000000000000",
962 => "000000000000000000000000",
963 => "000000000000000000000000",
964 => "000000000000000000000000",
965 => "000000000000000000000000",
966 => "000000000000000000000000",
967 => "000000000000000000000000",
968 => "000000000000000000000000",
969 => "000000000000000000000000",
970 => "000000000000000000000000",
971 => "000000000000000000000000",
972 => "000000000000000000000000",
973 => "000000000000000000000000",
974 => "000000000000000000000000",
975 => "000000000000000000000000",
976 => "000000000000000000000000",
977 => "000000000000000000000000",
978 => "000000000000000000000000",
979 => "000000000000000000000000",
980 => "000000000000000000000000",
981 => "000000000000000000000000",
982 => "000000000000000000000000",
983 => "000000000000000000000000",
984 => "000000000000000000000000",
985 => "000000000000000000000000",
986 => "000000000000000000000000",
987 => "000000000000000000000000",
988 => "000000000000000000000000",
989 => "000000000000000000000000",
990 => "000000000000000000000000",
991 => "000000000000000000000000",
992 => "000000000000000000000000",
993 => "000000000000000000000000",
994 => "000000000000000000000000",
995 => "000000000000000000000000",
996 => "000000000000000000000000",
997 => "000000000000000000000000",
998 => "000000000000000000000000",
999 => "000000000000000000000000",
1000 => "000000000000000000000000",
1001 => "000000000000000000000000",
1002 => "000000000000000000000000",
1003 => "000000000000000000000000",
1004 => "000000000000000000000000",
1005 => "000000000000000000000000",
1006 => "000000000000000000000000",
1007 => "000000000000000000000000",
1008 => "000000000000000000000000",
1009 => "000000000000000000000000",
1010 => "000000000000000000000000",
1011 => "000000000000000000000000",
1012 => "000000000000000000000000",
1013 => "000000000000000000000000",
1014 => "000000000000000000000000",
1015 => "000000000000000000000000",
1016 => "000000000000000000000000",
1017 => "000000000000000000000000",
1018 => "000000000000000000000000",
1019 => "000000000000000000000000",
1020 => "000000000000000000000000",
1021 => "000000000000000000000000",
1022 => "000000000000000000000000",
1023 => "000000000000000000000000",
1024 => "000000000000000000000000",
1025 => "000000000000000000000000",
1026 => "000000000000000000000000",
1027 => "000000000000000000000000",
1028 => "000000000000000000000000",
1029 => "000000000000000000000000",
1030 => "000000000000000000000000",
1031 => "000000000000000000000000",
1032 => "000000000000000000000000",
1033 => "000000000000000000000000",
1034 => "000000000000000000000000",
1035 => "000000000000000000000000",
1036 => "000000000000000000000000",
1037 => "000000000000000000000000",
1038 => "000000000000000000000000",
1039 => "000000000000000000000000",
1040 => "000000000000000000000000",
1041 => "000000000000000000000000",
1042 => "000000000000000000000000",
1043 => "000000000000000000000000",
1044 => "000000000000000000000000",
1045 => "000000000000000000000000",
1046 => "000000000000000000000000",
1047 => "000000000000000000000000",
1048 => "000000000000000000000000",
1049 => "000000000000000000000000",
1050 => "000000000000000000000000",
1051 => "000000000000000000000000",
1052 => "000000000000000000000000",
1053 => "000000000000000000000000",
1054 => "000000000000000000000000",
1055 => "000000000000000000000000",
1056 => "000000000000000000000000",
1057 => "000000000000000000000000",
1058 => "000000000000000000000000",
1059 => "000000000000000000000000",
1060 => "000000000000000000000000",
1061 => "000000000000000000000000",
1062 => "000000000000000000000000",
1063 => "000000000000000000000000",
1064 => "000000000000000000000000",
1065 => "000000000000000000000000",
1066 => "000000000000000000000000",
1067 => "000000000000000000000000",
1068 => "000000000000000000000000",
1069 => "000000000000000000000000",
1070 => "000000000000000000000000",
1071 => "000000000000000000000000",
1072 => "000000000000000000000000",
1073 => "000000000000000000000000",
1074 => "000000000000000000000000",
1075 => "000000000000000000000000",
1076 => "000000000000000000000000",
1077 => "000000000000000000000000",
1078 => "000000000000000000000000",
1079 => "000000000000000000000000",
1080 => "000000000000000000000000",
1081 => "000000000000000000000000",
1082 => "000000000000000000000000",
1083 => "000000000000000000000000",
1084 => "000000000000000000000000",
1085 => "000000000000000000000000",
1086 => "000000000000000000000000",
1087 => "000000000000000000000000",
1088 => "000000000000000000000000",
1089 => "000000000000000000000000",
1090 => "000000000000000000000000",
1091 => "000000000000000000000000",
1092 => "000000000000000000000000",
1093 => "000000000000000000000000",
1094 => "000000000000000000000000",
1095 => "000000000000000000000000",
1096 => "000000000000000000000000",
1097 => "000000000000000000000000",
1098 => "000000000000000000000000",
1099 => "000000000000000000000000",
1100 => "000000000000000000000000",
1101 => "000000000000000000000000",
1102 => "000000000000000000000000",
1103 => "000000000000000000000000",
1104 => "000000000000000000000000",
1105 => "000000000000000000000000",
1106 => "000000000000000000000000",
1107 => "000000000000000000000000",
1108 => "000000000000000000000000",
1109 => "000000000000000000000000",
1110 => "000000000000000000000000",
1111 => "000000000000000000000000",
1112 => "000000000000000000000000",
1113 => "000000000000000000000000",
1114 => "000000000000000000000000",
1115 => "000000000000000000000000",
1116 => "000000000000000000000000",
1117 => "000000000000000000000000",
1118 => "000000000000000000000000",
1119 => "000000000000000000000000",
1120 => "000000000000000000000000",
1121 => "000000000000000000000000",
1122 => "000000000000000000000000",
1123 => "000000000000000000000000",
1124 => "000000000000000000000000",
1125 => "000000000000000000000000",
1126 => "000000000000000000000000",
1127 => "000000000000000000000000",
1128 => "000000000000000000000000",
1129 => "000000000000000000000000",
1130 => "000000000000000000000000",
1131 => "000000000000000000000000",
1132 => "000000000000000000000000",
1133 => "000000000000000000000000",
1134 => "000000000000000000000000",
1135 => "000000000000000000000000",
1136 => "000000000000000000000000",
1137 => "000000000000000000000000",
1138 => "000000000000000000000000",
1139 => "000000000000000000000000",
1140 => "000000000000000000000000",
1141 => "000000000000000000000000",
1142 => "000000000000000000000000",
1143 => "000000000000000000000000",
1144 => "000000000000000000000000",
1145 => "000000000000000000000000",
1146 => "000000000000000000000000",
1147 => "000000000000000000000000",
1148 => "000000000000000000000000",
1149 => "000000000000000000000000",
1150 => "000000000000000000000000",
1151 => "000000000000000000000000",
1152 => "000000000000000000000000",
1153 => "000000000000000000000000",
1154 => "000000000000000000000000",
1155 => "000000000000000000000000",
1156 => "000000000000000000000000",
1157 => "000000000000000000000000",
1158 => "000000000000000000000000",
1159 => "000000000000000000000000",
1160 => "000000000000000000000000",
1161 => "000000000000000000000000",
1162 => "000000000000000000000000",
1163 => "000000000000000000000000",
1164 => "000000000000000000000000",
1165 => "000000000000000000000000",
1166 => "000000000000000000000000",
1167 => "000000000000000000000000",
1168 => "000000000000000000000000",
1169 => "000000000000000000000000",
1170 => "000000000000000000000000",
1171 => "000000000000000000000000",
1172 => "000000000000000000000000",
1173 => "000000000000000000000000",
1174 => "000000000000000000000000",
1175 => "000000000000000000000000",
1176 => "000000000000000000000000",
1177 => "000000000000000000000000",
1178 => "000000000000000000000000",
1179 => "000000000000000000000000",
1180 => "000000000000000000000000",
1181 => "000000000000000000000000",
1182 => "000000000000000000000000",
1183 => "000000000000000000000000",
1184 => "000000000000000000000000",
1185 => "000000000000000000000000",
1186 => "000000000000000000000000",
1187 => "000000000000000000000000",
1188 => "000000000000000000000000",
1189 => "000000000000000000000000",
1190 => "000000000000000000000000",
1191 => "000000000000000000000000",
1192 => "000000000000000000000000",
1193 => "000000000000000000000000",
1194 => "000000000000000000000000",
1195 => "000000000000000000000000",
1196 => "000000000000000000000000",
1197 => "000000000000000000000000",
1198 => "000000000000000000000000",
1199 => "000000000000000000000000",
1200 => "000000000000000000000000",
1201 => "000000000000000000000000",
1202 => "000000000000000000000000",
1203 => "000000000000000000000000",
1204 => "000000000000000000000000",
1205 => "000000000000000000000000",
1206 => "000000000000000000000000",
1207 => "000000000000000000000000",
1208 => "000000000000000000000000",
1209 => "000000000000000000000000",
1210 => "000000000000000000000000",
1211 => "000000000000000000000000",
1212 => "000000000000000000000000",
1213 => "000000000000000000000000",
1214 => "000000000000000000000000",
1215 => "000000000000000000000000",
1216 => "000000000000000000000000",
1217 => "000000000000000000000000",
1218 => "000000000000000000000000",
1219 => "000000000000000000000000",
1220 => "000000000000000000000000",
1221 => "000000000000000000000000",
1222 => "000000000000000000000000",
1223 => "000000000000000000000000",
1224 => "000000000000000000000000",
1225 => "000000000000000000000000",
1226 => "000000000000000000000000",
1227 => "000000000000000000000000",
1228 => "000000000000000000000000",
1229 => "000000000000000000000000",
1230 => "000000000000000000000000",
1231 => "000000000000000000000000",
1232 => "000000000000000000000000",
1233 => "000000000000000000000000",
1234 => "000000000000000000000000",
1235 => "000000000000000000000000",
1236 => "000000000000000000000000",
1237 => "000000000000000000000000",
1238 => "000000000000000000000000",
1239 => "000000000000000000000000",
1240 => "000000000000000000000000",
1241 => "000000000000000000000000",
1242 => "000000000000000000000000",
1243 => "000000000000000000000000",
1244 => "000000000000000000000000",
1245 => "000000000000000000000000",
1246 => "000000000000000000000000",
1247 => "000000000000000000000000",
1248 => "000000000000000000000000",
1249 => "000000000000000000000000",
1250 => "000000000000000000000000",
1251 => "000000000000000000000000",
1252 => "000000000000000000000000",
1253 => "000000000000000000000000",
1254 => "000000000000000000000000",
1255 => "000000000000000000000000",
1256 => "000000000000000000000000",
1257 => "000000000000000000000000",
1258 => "000000000000000000000000",
1259 => "000000000000000000000000",
1260 => "000000000000000000000000",
1261 => "000000000000000000000000",
1262 => "000000000000000000000000",
1263 => "000000000000000000000000",
1264 => "000000000000000000000000",
1265 => "000000000000000000000000",
1266 => "000000000000000000000000",
1267 => "000000000000000000000000",
1268 => "000000000000000000000000",
1269 => "000000000000000000000000",
1270 => "000000000000000000000000",
1271 => "000000000000000000000000",
1272 => "000000000000000000000000",
1273 => "000000000000000000000000",
1274 => "000000000000000000000000",
1275 => "000000000000000000000000",
1276 => "000000000000000000000000",
1277 => "000000000000000000000000",
1278 => "000000000000000000000000",
1279 => "000000000000000000000000",
1280 => "000000000000000000000000",
1281 => "000000000000000000000000",
1282 => "000000000000000000000000",
1283 => "000000000000000000000000",
1284 => "000000000000000000000000",
1285 => "000000000000000000000000",
1286 => "000000000000000000000000",
1287 => "000000000000000000000000",
1288 => "000000000000000000000000",
1289 => "000000000000000000000000",
1290 => "000000000000000000000000",
1291 => "000000000000000000000000",
1292 => "000000000000000000000000",
1293 => "000000000000000000000000",
1294 => "000000000000000000000000",
1295 => "000000000000000000000000",
1296 => "000000000000000000000000",
1297 => "000000000000000000000000",
1298 => "000000000000000000000000",
1299 => "000000000000000000000000",
1300 => "000000000000000000000000",
1301 => "000000000000000000000000",
1302 => "000000000000000000000000",
1303 => "000000000000000000000000",
1304 => "000000000000000000000000",
1305 => "000000000000000000000000",
1306 => "000000000000000000000000",
1307 => "000000000000000000000000",
1308 => "000000000000000000000000",
1309 => "000000000000000000000000",
1310 => "000000000000000000000000",
1311 => "000000000000000000000000",
1312 => "000000000000000000000000",
1313 => "000000000000000000000000",
1314 => "000000000000000000000000",
1315 => "000000000000000000000000",
1316 => "000000000000000000000000",
1317 => "000000000000000000000000",
1318 => "000000000000000000000000",
1319 => "000000000000000000000000",
1320 => "000000000000000000000000",
1321 => "000000000000000000000000",
1322 => "000000000000000000000000",
1323 => "000000000000000000000000",
1324 => "000000000000000000000000",
1325 => "000000000000000000000000",
1326 => "000000000000000000000000",
1327 => "000000000000000000000000",
1328 => "000000000000000000000000",
1329 => "000000000000000000000000",
1330 => "000000000000000000000000",
1331 => "000000000000000000000000",
1332 => "000000000000000000000000",
1333 => "000000000000000000000000",
1334 => "000000000000000000000000",
1335 => "000000000000000000000000",
1336 => "000000000000000000000000",
1337 => "000000000000000000000000",
1338 => "000000000000000000000000",
1339 => "000000000000000000000000",
1340 => "000000000000000000000000",
1341 => "000000000000000000000000",
1342 => "000000000000000000000000",
1343 => "000000000000000000000000",
1344 => "000000000000000000000000",
1345 => "000000000000000000000000",
1346 => "000000000000000000000000",
1347 => "000000000000000000000000",
1348 => "000000000000000000000000",
1349 => "000000000000000000000000",
1350 => "000000000000000000000000",
1351 => "000000000000000000000000",
1352 => "000000000000000000000000",
1353 => "000000000000000000000000",
1354 => "000000000000000000000000",
1355 => "000000000000000000000000",
1356 => "000000000000000000000000",
1357 => "000000000000000000000000",
1358 => "000000000000000000000000",
1359 => "000000000000000000000000",
1360 => "000000000000000000000000",
1361 => "000000000000000000000000",
1362 => "000000000000000000000000",
1363 => "000000000000000000000000",
1364 => "000000000000000000000000",
1365 => "000000000000000000000000",
1366 => "000000000000000000000000",
1367 => "000000000000000000000000",
1368 => "000000000000000000000000",
1369 => "000000000000000000000000",
1370 => "000000000000000000000000",
1371 => "000000000000000000000000",
1372 => "000000000000000000000000",
1373 => "000000000000000000000000",
1374 => "000000000000000000000000",
1375 => "000000000000000000000000",
1376 => "000000000000000000000000",
1377 => "000000000000000000000000",
1378 => "000000000000000000000000",
1379 => "000000000000000000000000",
1380 => "000000000000000000000000",
1381 => "000000000000000000000000",
1382 => "000000000000000000000000",
1383 => "000000000000000000000000",
1384 => "000000000000000000000000",
1385 => "000000000000000000000000",
1386 => "000000000000000000000000",
1387 => "000000000000000000000000",
1388 => "000000000000000000000000",
1389 => "000000000000000000000000",
1390 => "000000000000000000000000",
1391 => "000000000000000000000000",
1392 => "000000000000000000000000",
1393 => "000000000000000000000000",
1394 => "000000000000000000000000",
1395 => "000000000000000000000000",
1396 => "000000000000000000000000",
1397 => "000000000000000000000000",
1398 => "000000000000000000000000",
1399 => "000000000000000000000000",
1400 => "000000000000000000000000",
1401 => "000000000000000000000000",
1402 => "000000000000000000000000",
1403 => "000000000000000000000000",
1404 => "000000000000000000000000",
1405 => "000000000000000000000000",
1406 => "000000000000000000000000",
1407 => "000000000000000000000000",
1408 => "000000000000000000000000",
1409 => "000000000000000000000000",
1410 => "000000000000000000000000",
1411 => "000000000000000000000000",
1412 => "000000000000000000000000",
1413 => "000000000000000000000000",
1414 => "000000000000000000000000",
1415 => "000000000000000000000000",
1416 => "000000000000000000000000",
1417 => "000000000000000000000000",
1418 => "000000000000000000000000",
1419 => "000000000000000000000000",
1420 => "000000000000000000000000",
1421 => "000000000000000000000000",
1422 => "000000000000000000000000",
1423 => "000000000000000000000000",
1424 => "000000000000000000000000",
1425 => "000000000000000000000000",
1426 => "000000000000000000000000",
1427 => "000000000000000000000000",
1428 => "000000000000000000000000",
1429 => "000000000000000000000000",
1430 => "000000000000000000000000",
1431 => "000000000000000000000000",
1432 => "000000000000000000000000",
1433 => "000000000000000000000000",
1434 => "000000000000000000000000",
1435 => "000000000000000000000000",
1436 => "000000000000000000000000",
1437 => "000000000000000000000000",
1438 => "000000000000000000000000",
1439 => "000000000000000000000000",
1440 => "000000000000000000000000",
1441 => "000000000000000000000000",
1442 => "000000000000000000000000",
1443 => "000000000000000000000000",
1444 => "000000000000000000000000",
1445 => "000000000000000000000000",
1446 => "000000000000000000000000",
1447 => "000000000000000000000000",
1448 => "000000000000000000000000",
1449 => "000000000000000000000000",
1450 => "000000000000000000000000",
1451 => "000000000000000000000000",
1452 => "000000000000000000000000",
1453 => "000000000000000000000000",
1454 => "000000000000000000000000",
1455 => "000000000000000000000000",
1456 => "000000000000000000000000",
1457 => "000000000000000000000000",
1458 => "000000000000000000000000",
1459 => "000000000000000000000000",
1460 => "000000000000000000000000",
1461 => "000000000000000000000000",
1462 => "000000000000000000000000",
1463 => "000000000000000000000000",
1464 => "000000000000000000000000",
1465 => "000000000000000000000000",
1466 => "000000000000000000000000",
1467 => "000000000000000000000000",
1468 => "000000000000000000000000",
1469 => "000000000000000000000000",
1470 => "000000000000000000000000",
1471 => "000000000000000000000000",
1472 => "000000000000000000000000",
1473 => "000000000000000000000000",
1474 => "000000000000000000000000",
1475 => "000000000000000000000000",
1476 => "000000000000000000000000",
1477 => "000000000000000000000000",
1478 => "000000000000000000000000",
1479 => "000000000000000000000000",
1480 => "000000000000000000000000",
1481 => "000000000000000000000000",
1482 => "000000000000000000000000",
1483 => "000000000000000000000000",
1484 => "000000000000000000000000",
1485 => "000000000000000000000000",
1486 => "000000000000000000000000",
1487 => "000000000000000000000000",
1488 => "000000000000000000000000",
1489 => "000000000000000000000000",
1490 => "000000000000000000000000",
1491 => "000000000000000000000000",
1492 => "000000000000000000000000",
1493 => "000000000000000000000000",
1494 => "000000000000000000000000",
1495 => "000000000000000000000000",
1496 => "000000000000000000000000",
1497 => "000000000000000000000000",
1498 => "000000000000000000000000",
1499 => "000000000000000000000000",
1500 => "000000000000000000000000",
1501 => "000000000000000000000000",
1502 => "000000000000000000000000",
1503 => "000000000000000000000000",
1504 => "000000000000000000000000",
1505 => "000000000000000000000000",
1506 => "000000000000000000000000",
1507 => "000000000000000000000000",
1508 => "000000000000000000000000",
1509 => "000000000000000000000000",
1510 => "000000000000000000000000",
1511 => "000000000000000000000000",
1512 => "000000000000000000000000",
1513 => "000000000000000000000000",
1514 => "000000000000000000000000",
1515 => "000000000000000000000000",
1516 => "000000000000000000000000",
1517 => "000000000000000000000000",
1518 => "000000000000000000000000",
1519 => "000000000000000000000000",
1520 => "000000000000000000000000",
1521 => "000000000000000000000000",
1522 => "000000000000000000000000",
1523 => "000000000000000000000000",
1524 => "000000000000000000000000",
1525 => "000000000000000000000000",
1526 => "000000000000000000000000",
1527 => "000000000000000000000000",
1528 => "000000000000000000000000",
1529 => "000000000000000000000000",
1530 => "000000000000000000000000",
1531 => "000000000000000000000000",
1532 => "000000000000000000000000",
1533 => "000000000000000000000000",
1534 => "000000000000000000000000",
1535 => "000000000000000000000000",
1536 => "000000000000000000000000",
1537 => "000000000000000000000000",
1538 => "000000000000000000000000",
1539 => "000000000000000000000000",
1540 => "000000000000000000000000",
1541 => "000000000000000000000000",
1542 => "000000000000000000000000",
1543 => "000000000000000000000000",
1544 => "000000000000000000000000",
1545 => "000000000000000000000000",
1546 => "000000000000000000000000",
1547 => "000000000000000000000000",
1548 => "000000000000000000000000",
1549 => "000000000000000000000000",
1550 => "000000000000000000000000",
1551 => "000000000000000000000000",
1552 => "000000000000000000000000",
1553 => "000000000000000000000000",
1554 => "000000000000000000000000",
1555 => "000000000000000000000000",
1556 => "000000000000000000000000",
1557 => "000000000000000000000000",
1558 => "000000000000000000000000",
1559 => "000000000000000000000000",
1560 => "000000000000000000000000",
1561 => "000000000000000000000000",
1562 => "000000000000000000000000",
1563 => "000000000000000000000000",
1564 => "000000000000000000000000",
1565 => "000000000000000000000000",
1566 => "000000000000000000000000",
1567 => "000000000000000000000000",
1568 => "000000000000000000000000",
1569 => "000000000000000000000000",
1570 => "000000000000000000000000",
1571 => "000000000000000000000000",
1572 => "000000000000000000000000",
1573 => "000000000000000000000000",
1574 => "000000000000000000000000",
1575 => "000000000000000000000000",
1576 => "000000000000000000000000",
1577 => "000000000000000000000000",
1578 => "000000000000000000000000",
1579 => "000000000000000000000000",
1580 => "000000000000000000000000",
1581 => "000000000000000000000000",
1582 => "000000000000000000000000",
1583 => "000000000000000000000000",
1584 => "000000000000000000000000",
1585 => "000000000000000000000000",
1586 => "000000000000000000000000",
1587 => "000000000000000000000000",
1588 => "000000000000000000000000",
1589 => "000000000000000000000000",
1590 => "000000000000000000000000",
1591 => "000000000000000000000000",
1592 => "000000000000000000000000",
1593 => "000000000000000000000000",
1594 => "000000000000000000000000",
1595 => "000000000000000000000000",
1596 => "000000000000000000000000",
1597 => "000000000000000000000000",
1598 => "000000000000000000000000",
1599 => "000000000000000000000000",
1600 => "000000000000000000000000",
1601 => "000000000000000000000000",
1602 => "000000000000000000000000",
1603 => "000000000000000000000000",
1604 => "000000000000000000000000",
1605 => "000000000000000000000000",
1606 => "000000000000000000000000",
1607 => "000000000000000000000000",
1608 => "000000000000000000000000",
1609 => "000000000000000000000000",
1610 => "000000000000000000000000",
1611 => "000000000000000000000000",
1612 => "000000000000000000000000",
1613 => "000000000000000000000000",
1614 => "000000000000000000000000",
1615 => "000000000000000000000000",
1616 => "000000000000000000000000",
1617 => "000000000000000000000000",
1618 => "000000000000000000000000",
1619 => "000000000000000000000000",
1620 => "000000000000000000000000",
1621 => "000000000000000000000000",
1622 => "000000000000000000000000",
1623 => "000000000000000000000000",
1624 => "000000000000000000000000",
1625 => "000000000000000000000000",
1626 => "000000000000000000000000",
1627 => "000000000000000000000000",
1628 => "000000000000000000000000",
1629 => "000000000000000000000000",
1630 => "000000000000000000000000",
1631 => "000000000000000000000000",
1632 => "000000000000000000000000",
1633 => "000000000000000000000000",
1634 => "000000000000000000000000",
1635 => "000000000000000000000000",
1636 => "000000000000000000000000",
1637 => "000000000000000000000000",
1638 => "000000000000000000000000",
1639 => "000000000000000000000000",
1640 => "000000000000000000000000",
1641 => "000000000000000000000000",
1642 => "000000000000000000000000",
1643 => "000000000000000000000000",
1644 => "000000000000000000000000",
1645 => "000000000000000000000000",
1646 => "000000000000000000000000",
1647 => "000000000000000000000000",
1648 => "000000000000000000000000",
1649 => "000000000000000000000000",
1650 => "000000000000000000000000",
1651 => "000000000000000000000000",
1652 => "000000000000000000000000",
1653 => "000000000000000000000000",
1654 => "000000000000000000000000",
1655 => "000000000000000000000000",
1656 => "000000000000000000000000",
1657 => "000000000000000000000000",
1658 => "000000000000000000000000",
1659 => "000000000000000000000000",
1660 => "000000000000000000000000",
1661 => "000000000000000000000000",
1662 => "000000000000000000000000",
1663 => "000000000000000000000000",
1664 => "000000000000000000000000",
1665 => "000000000000000000000000",
1666 => "000000000000000000000000",
1667 => "000000000000000000000000",
1668 => "000000000000000000000000",
1669 => "000000000000000000000000",
1670 => "000000000000000000000000",
1671 => "000000000000000000000000",
1672 => "000000000000000000000000",
1673 => "000000000000000000000000",
1674 => "000000000000000000000000",
1675 => "000000000000000000000000",
1676 => "000000000000000000000000",
1677 => "000000000000000000000000",
1678 => "000000000000000000000000",
1679 => "000000000000000000000000",
1680 => "000000000000000000000000",
1681 => "000000000000000000000000",
1682 => "000000000000000000000000",
1683 => "000000000000000000000000",
1684 => "000000000000000000000000",
1685 => "000000000000000000000000",
1686 => "000000000000000000000000",
1687 => "000000000000000000000000",
1688 => "000000000000000000000000",
1689 => "000000000000000000000000",
1690 => "000000000000000000000000",
1691 => "000000000000000000000000",
1692 => "000000000000000000000000",
1693 => "000000000000000000000000",
1694 => "000000000000000000000000",
1695 => "000000000000000000000000",
1696 => "000000000000000000000000",
1697 => "000000000000000000000000",
1698 => "000000000000000000000000",
1699 => "000000000000000000000000",
1700 => "000000000000000000000000",
1701 => "000000000000000000000000",
1702 => "000000000000000000000000",
1703 => "000000000000000000000000",
1704 => "000000000000000000000000",
1705 => "000000000000000000000000",
1706 => "000000000000000000000000",
1707 => "000000000000000000000000",
1708 => "000000000000000000000000",
1709 => "000000000000000000000000",
1710 => "000000000000000000000000",
1711 => "000000000000000000000000",
1712 => "000000000000000000000000",
1713 => "000000000000000000000000",
1714 => "000000000000000000000000",
1715 => "000000000000000000000000",
1716 => "000000000000000000000000",
1717 => "000000000000000000000000",
1718 => "000000000000000000000000",
1719 => "000000000000000000000000",
1720 => "000000000000000000000000",
1721 => "000000000000000000000000",
1722 => "000000000000000000000000",
1723 => "000000000000000000000000",
1724 => "000000000000000000000000",
1725 => "000000000000000000000000",
1726 => "000000000000000000000000",
1727 => "000000000000000000000000",
1728 => "000000000000000000000000",
1729 => "000000000000000000000000",
1730 => "000000000000000000000000",
1731 => "000000000000000000000000",
1732 => "000000000000000000000000",
1733 => "000000000000000000000000",
1734 => "000000000000000000000000",
1735 => "000000000000000000000000",
1736 => "000000000000000000000000",
1737 => "000000000000000000000000",
1738 => "000000000000000000000000",
1739 => "000000000000000000000000",
1740 => "000000000000000000000000",
1741 => "000000000000000000000000",
1742 => "000000000000000000000000",
1743 => "000000000000000000000000",
1744 => "000000000000000000000000",
1745 => "000000000000000000000000",
1746 => "000000000000000000000000",
1747 => "000000000000000000000000",
1748 => "000000000000000000000000",
1749 => "000000000000000000000000",
1750 => "000000000000000000000000",
1751 => "000000000000000000000000",
1752 => "000000000000000000000000",
1753 => "000000000000000000000000",
1754 => "000000000000000000000000",
1755 => "000000000000000000000000",
1756 => "000000000000000000000000",
1757 => "000000000000000000000000",
1758 => "000000000000000000000000",
1759 => "000000000000000000000000",
1760 => "000000000000000000000000",
1761 => "000000000000000000000000",
1762 => "000000000000000000000000",
1763 => "000000000000000000000000",
1764 => "000000000000000000000000",
1765 => "000000000000000000000000",
1766 => "000000000000000000000000",
1767 => "000000000000000000000000",
1768 => "000000000000000000000000",
1769 => "000000000000000000000000",
1770 => "000000000000000000000000",
1771 => "000000000000000000000000",
1772 => "000000000000000000000000",
1773 => "000000000000000000000000",
1774 => "000000000000000000000000",
1775 => "000000000000000000000000",
1776 => "000000000000000000000000",
1777 => "000000000000000000000000",
1778 => "000000000000000000000000",
1779 => "000000000000000000000000",
1780 => "000000000000000000000000",
1781 => "000000000000000000000000",
1782 => "000000000000000000000000",
1783 => "000000000000000000000000",
1784 => "000000000000000000000000",
1785 => "000000000000000000000000",
1786 => "000000000000000000000000",
1787 => "000000000000000000000000",
1788 => "000000000000000000000000",
1789 => "000000000000000000000000",
1790 => "000000000000000000000000",
1791 => "000000000000000000000000",
1792 => "000000000000000000000000",
1793 => "000000000000000000000000",
1794 => "000000000000000000000000",
1795 => "000000000000000000000000",
1796 => "000000000000000000000000",
1797 => "000000000000000000000000",
1798 => "000000000000000000000000",
1799 => "000000000000000000000000",
1800 => "000000000000000000000000",
1801 => "000000000000000000000000",
1802 => "000000000000000000000000",
1803 => "000000000000000000000000",
1804 => "000000000000000000000000",
1805 => "000000000000000000000000",
1806 => "000000000000000000000000",
1807 => "000000000000000000000000",
1808 => "000000000000000000000000",
1809 => "000000000000000000000000",
1810 => "000000000000000000000000",
1811 => "000000000000000000000000",
1812 => "000000000000000000000000",
1813 => "000000000000000000000000",
1814 => "000000000000000000000000",
1815 => "000000000000000000000000",
1816 => "000000000000000000000000",
1817 => "000000000000000000000000",
1818 => "000000000000000000000000",
1819 => "000000000000000000000000",
1820 => "000000000000000000000000",
1821 => "000000000000000000000000",
1822 => "000000000000000000000000",
1823 => "000000000000000000000000",
1824 => "000000000000000000000000",
1825 => "000000000000000000000000",
1826 => "000000000000000000000000",
1827 => "000000000000000000000000",
1828 => "000000000000000000000000",
1829 => "000000000000000000000000",
1830 => "000000000000000000000000",
1831 => "000000000000000000000000",
1832 => "000000000000000000000000",
1833 => "000000000000000000000000",
1834 => "000000000000000000000000",
1835 => "000000000000000000000000",
1836 => "000000000000000000000000",
1837 => "000000000000000000000000",
1838 => "000000000000000000000000",
1839 => "000000000000000000000000",
1840 => "000000000000000000000000",
1841 => "000000000000000000000000",
1842 => "000000000000000000000000",
1843 => "000000000000000000000000",
1844 => "000000000000000000000000",
1845 => "000000000000000000000000",
1846 => "000000000000000000000000",
1847 => "000000000000000000000000",
1848 => "000000000000000000000000",
1849 => "000000000000000000000000",
1850 => "000000000000000000000000",
1851 => "000000000000000000000000",
1852 => "000000000000000000000000",
1853 => "000000000000000000000000",
1854 => "000000000000000000000000",
1855 => "000000000000000000000000",
1856 => "000000000000000000000000",
1857 => "000000000000000000000000",
1858 => "000000000000000000000000",
1859 => "000000000000000000000000",
1860 => "000000000000000000000000",
1861 => "000000000000000000000000",
1862 => "000000000000000000000000",
1863 => "000000000000000000000000",
1864 => "000000000000000000000000",
1865 => "000000000000000000000000",
1866 => "000000000000000000000000",
1867 => "000000000000000000000000",
1868 => "000000000000000000000000",
1869 => "000000000000000000000000",
1870 => "000000000000000000000000",
1871 => "000000000000000000000000",
1872 => "000000000000000000000000",
1873 => "000000000000000000000000",
1874 => "000000000000000000000000",
1875 => "000000000000000000000000",
1876 => "000000000000000000000000",
1877 => "000000000000000000000000",
1878 => "000000000000000000000000",
1879 => "000000000000000000000000",
1880 => "000000000000000000000000",
1881 => "000000000000000000000000",
1882 => "000000000000000000000000",
1883 => "000000000000000000000000",
1884 => "000000000000000000000000",
1885 => "000000000000000000000000",
1886 => "000000000000000000000000",
1887 => "000000000000000000000000",
1888 => "000000000000000000000000",
1889 => "000000000000000000000000",
1890 => "000000000000000000000000",
1891 => "000000000000000000000000",
1892 => "000000000000000000000000",
1893 => "000000000000000000000000",
1894 => "000000000000000000000000",
1895 => "000000000000000000000000",
1896 => "000000000000000000000000",
1897 => "000000000000000000000000",
1898 => "000000000000000000000000",
1899 => "000000000000000000000000",
1900 => "000000000000000000000000",
1901 => "000000000000000000000000",
1902 => "000000000000000000000000",
1903 => "000000000000000000000000",
1904 => "000000000000000000000000",
1905 => "000000000000000000000000",
1906 => "000000000000000000000000",
1907 => "000000000000000000000000",
1908 => "000000000000000000000000",
1909 => "000000000000000000000000",
1910 => "000000000000000000000000",
1911 => "000000000000000000000000",
1912 => "000000000000000000000000",
1913 => "000000000000000000000000",
1914 => "000000000000000000000000",
1915 => "000000000000000000000000",
1916 => "000000000000000000000000",
1917 => "000000000000000000000000",
1918 => "000000000000000000000000",
1919 => "000000000000000000000000",
1920 => "000000000000000000000000",
1921 => "000000000000000000000000",
1922 => "000000000000000000000000",
1923 => "000000000000000000000000",
1924 => "000000000000000000000000",
1925 => "000000000000000000000000",
1926 => "000000000000000000000000",
1927 => "000000000000000000000000",
1928 => "000000000000000000000000",
1929 => "000000000000000000000000",
1930 => "000000000000000000000000",
1931 => "000000000000000000000000",
1932 => "000000000000000000000000",
1933 => "000000000000000000000000",
1934 => "000000000000000000000000",
1935 => "000000000000000000000000",
1936 => "000000000000000000000000",
1937 => "000000000000000000000000",
1938 => "000000000000000000000000",
1939 => "000000000000000000000000",
1940 => "000000000000000000000000",
1941 => "000000000000000000000000",
1942 => "000000000000000000000000",
1943 => "000000000000000000000000",
1944 => "000000000000000000000000",
1945 => "000000000000000000000000",
1946 => "000000000000000000000000",
1947 => "000000000000000000000000",
1948 => "000000000000000000000000",
1949 => "000000000000000000000000",
1950 => "000000000000000000000000",
1951 => "000000000000000000000000",
1952 => "000000000000000000000000",
1953 => "000000000000000000000000",
1954 => "000000000000000000000000",
1955 => "000000000000000000000000",
1956 => "000000000000000000000000",
1957 => "000000000000000000000000",
1958 => "000000000000000000000000",
1959 => "000000000000000000000000",
1960 => "000000000000000000000000",
1961 => "000000000000000000000000",
1962 => "000000000000000000000000",
1963 => "000000000000000000000000",
1964 => "000000000000000000000000",
1965 => "000000000000000000000000",
1966 => "000000000000000000000000",
1967 => "000000000000000000000000",
1968 => "000000000000000000000000",
1969 => "000000000000000000000000",
1970 => "000000000000000000000000",
1971 => "000000000000000000000000",
1972 => "000000000000000000000000",
1973 => "000000000000000000000000",
1974 => "000000000000000000000000",
1975 => "000000000000000000000000",
1976 => "000000000000000000000000",
1977 => "000000000000000000000000",
1978 => "000000000000000000000000",
1979 => "000000000000000000000000",
1980 => "000000000000000000000000",
1981 => "000000000000000000000000",
1982 => "000000000000000000000000",
1983 => "000000000000000000000000",
1984 => "000000000000000000000000",
1985 => "000000000000000000000000",
1986 => "000000000000000000000000",
1987 => "000000000000000000000000",
1988 => "000000000000000000000000",
1989 => "000000000000000000000000",
1990 => "000000000000000000000000",
1991 => "000000000000000000000000",
1992 => "000000000000000000000000",
1993 => "000000000000000000000000",
1994 => "000000000000000000000000",
1995 => "000000000000000000000000",
1996 => "000000000000000000000000",
1997 => "000000000000000000000000",
1998 => "000000000000000000000000",
1999 => "000000000000000000000000",
2000 => "000000000000000000000000",
2001 => "000000000000000000000000",
2002 => "000000000000000000000000",
2003 => "000000000000000000000000",
2004 => "000000000000000000000000",
2005 => "000000000000000000000000",
2006 => "000000000000000000000000",
2007 => "000000000000000000000000",
2008 => "000000000000000000000000",
2009 => "000000000000000000000000",
2010 => "000000000000000000000000",
2011 => "000000000000000000000000",
2012 => "000000000000000000000000",
2013 => "000000000000000000000000",
2014 => "000000000000000000000000",
2015 => "000000000000000000000000",
2016 => "000000000000000000000000",
2017 => "000000000000000000000000",
2018 => "000000000000000000000000",
2019 => "000000000000000000000000",
2020 => "000000000000000000000000",
2021 => "000000000000000000000000",
2022 => "000000000000000000000000",
2023 => "000000000000000000000000",
2024 => "000000000000000000000000",
2025 => "000000000000000000000000",
2026 => "000000000000000000000000",
2027 => "000000000000000000000000",
2028 => "000000000000000000000000",
2029 => "000000000000000000000000",
2030 => "000000000000000000000000",
2031 => "000000000000000000000000",
2032 => "000000000000000000000000",
2033 => "000000000000000000000000",
2034 => "000000000000000000000000",
2035 => "000000000000000000000000",
2036 => "000000000000000000000000",
2037 => "000000000000000000000000",
2038 => "000000000000000000000000",
2039 => "000000000000000000000000",
2040 => "000000000000000000000000",
2041 => "000000000000000000000000",
2042 => "000000000000000000000000",
2043 => "000000000000000000000000",
2044 => "000000000000000000000000",
2045 => "000000000000000000000000",
2046 => "000000000000000000000000",
2047 => "000000000000000000000000",
2048 => "000000000000000000000000",
2049 => "000000000000000000000000",
2050 => "000000000000000000000000",
2051 => "000000000000000000000000",
2052 => "000000000000000000000000",
2053 => "000000000000000000000000",
2054 => "000000000000000000000000",
2055 => "000000000000000000000000",
2056 => "000000000000000000000000",
2057 => "000000000000000000000000",
2058 => "000000000000000000000000",
2059 => "000000000000000000000000",
2060 => "000000000000000000000000",
2061 => "000000000000000000000000",
2062 => "000000000000000000000000",
2063 => "000000000000000000000000",
2064 => "000000000000000000000000",
2065 => "000000000000000000000000",
2066 => "000000000000000000000000",
2067 => "000000000000000000000000",
2068 => "000000000000000000000000",
2069 => "000000000000000000000000",
2070 => "000000000000000000000000",
2071 => "000000000000000000000000",
2072 => "000000000000000000000000",
2073 => "000000000000000000000000",
2074 => "000000000000000000000000",
2075 => "000000000000000000000000",
2076 => "000000000000000000000000",
2077 => "000000000000000000000000",
2078 => "000000000000000000000000",
2079 => "000000000000000000000000",
2080 => "000000000000000000000000",
2081 => "000000000000000000000000",
2082 => "000000000000000000000000",
2083 => "000000000000000000000000",
2084 => "000000000000000000000000",
2085 => "000000000000000000000000",
2086 => "000000000000000000000000",
2087 => "000000000000000000000000",
2088 => "000000000000000000000000",
2089 => "000000000000000000000000",
2090 => "000000000000000000000000",
2091 => "000000000000000000000000",
2092 => "000000000000000000000000",
2093 => "000000000000000000000000",
2094 => "000000000000000000000000",
2095 => "000000000000000000000000",
2096 => "000000000000000000000000",
2097 => "000000000000000000000000",
2098 => "000000000000000000000000",
2099 => "000000000000000000000000",
2100 => "000000000000000000000000",
2101 => "000000000000000000000000",
2102 => "000000000000000000000000",
2103 => "000000000000000000000000",
2104 => "000000000000000000000000",
2105 => "000000000000000000000000",
2106 => "000000000000000000000000",
2107 => "000000000000000000000000",
2108 => "000000000000000000000000",
2109 => "000000000000000000000000",
2110 => "000000000000000000000000",
2111 => "000000000000000000000000",
2112 => "000000000000000000000000",
2113 => "000000000000000000000000",
2114 => "000000000000000000000000",
2115 => "000000000000000000000000",
2116 => "000000000000000000000000",
2117 => "000000000000000000000000",
2118 => "000000000000000000000000",
2119 => "000000000000000000000000",
2120 => "000000000000000000000000",
2121 => "000000000000000000000000",
2122 => "000000000000000000000000",
2123 => "000000000000000000000000",
2124 => "000000000000000000000000",
2125 => "000000000000000000000000",
2126 => "000000000000000000000000",
2127 => "000000000000000000000000",
2128 => "000000000000000000000000",
2129 => "000000000000000000000000",
2130 => "000000000000000000000000",
2131 => "000000000000000000000000",
2132 => "000000000000000000000000",
2133 => "000000000000000000000000",
2134 => "000000000000000000000000",
2135 => "000000000000000000000000",
2136 => "000000000000000000000000",
2137 => "000000000000000000000000",
2138 => "000000000000000000000000",
2139 => "000000000000000000000000",
2140 => "000000000000000000000000",
2141 => "000000000000000000000000",
2142 => "000000000000000000000000",
2143 => "000000000000000000000000",
2144 => "000000000000000000000000",
2145 => "000000000000000000000000",
2146 => "000000000000000000000000",
2147 => "000000000000000000000000",
2148 => "000000000000000000000000",
2149 => "000000000000000000000000",
2150 => "000000000000000000000000",
2151 => "000000000000000000000000",
2152 => "000000000000000000000000",
2153 => "000000000000000000000000",
2154 => "000000000000000000000000",
2155 => "000000000000000000000000",
2156 => "000000000000000000000000",
2157 => "000000000000000000000000",
2158 => "000000000000000000000000",
2159 => "000000000000000000000000",
2160 => "000000000000000000000000",
2161 => "000000000000000000000000",
2162 => "000000000000000000000000",
2163 => "000000000000000000000000",
2164 => "000000000000000000000000",
2165 => "000000000000000000000000",
2166 => "000000000000000000000000",
2167 => "000000100000001000000010",
2168 => "010000100100001001000010",
2169 => "010000100100001001000010",
2170 => "000101010001010100010101",
2171 => "000000000000000000000000",
2172 => "000000000000000000000000",
2173 => "000000000000000000000000",
2174 => "000000000000000000000000",
2175 => "000000000000000000000000",
2176 => "000000000000000000000000",
2177 => "000000000000000000000000",
2178 => "000000000000000000000000",
2179 => "000000000000000000000000",
2180 => "000000000000000000000000",
2181 => "000000000000000000000000",
2182 => "000000000000000000000000",
2183 => "000000000000000000000000",
2184 => "000000000000000000000000",
2185 => "000000000000000000000000",
2186 => "000000000000000000000000",
2187 => "000000000000000000000000",
2188 => "000000000000000000000000",
2189 => "000000000000000000000000",
2190 => "000000000000000000000000",
2191 => "000000000000000000000000",
2192 => "000000000000000000000000",
2193 => "000000000000000000000000",
2194 => "000000000000000000000000",
2195 => "000000000000000000000000",
2196 => "000000000000000000000000",
2197 => "000000000000000000000000",
2198 => "000000000000000000000000",
2199 => "000000000000000000000000",
2200 => "000000000000000000000000",
2201 => "000000000000000000000000",
2202 => "000000000000000000000000",
2203 => "000000000000000000000000",
2204 => "000000000000000000000000",
2205 => "000000000000000000000000",
2206 => "000000000000000000000000",
2207 => "000000000000000000000000",
2208 => "000000000000000000000000",
2209 => "000000000000000000000000",
2210 => "000000000000000000000000",
2211 => "000000000000000000000000",
2212 => "000000000000000000000000",
2213 => "000000000000000000000000",
2214 => "000000000000000000000000",
2215 => "000000000000000000000000",
2216 => "000000000000000000000000",
2217 => "000000000000000000000000",
2218 => "000000000000000000000000",
2219 => "000000000000000000000000",
2220 => "000000000000000000000000",
2221 => "000000000000000000000000",
2222 => "000000000000000000000000",
2223 => "000000000000000000000000",
2224 => "000000000000000000000000",
2225 => "000000000000000000000000",
2226 => "000000000000000000000000",
2227 => "000000000000000000000000",
2228 => "000000000000000000000000",
2229 => "000000000000000000000000",
2230 => "000000000000000000000000",
2231 => "000000000000000000000000",
2232 => "000000000000000000000000",
2233 => "000000000000000000000000",
2234 => "000000000000000000000000",
2235 => "000000000000000000000000",
2236 => "000000000000000000000000",
2237 => "000000000000000000000000",
2238 => "000000000000000000000000",
2239 => "000000000000000000000000",
2240 => "000000000000000000000000",
2241 => "000000000000000000000000",
2242 => "000000000000000000000000",
2243 => "000000000000000000000000",
2244 => "000000000000000000000000",
2245 => "000000000000000000000000",
2246 => "000000000000000000000000",
2247 => "000000000000000000000000",
2248 => "000000000000000000000000",
2249 => "000000000000000000000000",
2250 => "000000000000000000000000",
2251 => "000000000000000000000000",
2252 => "000000000000000000000000",
2253 => "000000000000000000000000",
2254 => "000000000000000000000000",
2255 => "000000000000000000000000",
2256 => "000000000000000000000000",
2257 => "000000000000000000000000",
2258 => "000000000000000000000000",
2259 => "000000000000000000000000",
2260 => "000000000000000000000000",
2261 => "000000000000000000000000",
2262 => "000000000000000000000000",
2263 => "000000000000000000000000",
2264 => "000000000000000000000000",
2265 => "000000000000000000000000",
2266 => "000000000000000000000000",
2267 => "000000000000000000000000",
2268 => "000000000000000000000000",
2269 => "000000000000000000000000",
2270 => "000000000000000000000000",
2271 => "000000000000000000000000",
2272 => "000000000000000000000000",
2273 => "000000000000000000000000",
2274 => "000000000000000000000000",
2275 => "000000000000000000000000",
2276 => "000000000000000000000000",
2277 => "000000000000000000000000",
2278 => "000000000000000000000000",
2279 => "000000000000000000000000",
2280 => "000000000000000000000000",
2281 => "000000000000000000000000",
2282 => "000000000000000000000000",
2283 => "000000000000000000000000",
2284 => "000000000000000000000000",
2285 => "000000000000000000000000",
2286 => "000000000000000000000000",
2287 => "000000000000000000000000",
2288 => "000000000000000000000000",
2289 => "000000000000000000000000",
2290 => "000000000000000000000000",
2291 => "000000000000000000000000",
2292 => "000000000000000000000000",
2293 => "000000000000000000000000",
2294 => "000000000000000000000000",
2295 => "000000000000000000000000",
2296 => "000000000000000000000000",
2297 => "000000000000000000000000",
2298 => "000000000000000000000000",
2299 => "000000000000000000000000",
2300 => "000000000000000000000000",
2301 => "000000000000000000000000",
2302 => "000000000000000000000000",
2303 => "000000000000000000000000",
2304 => "000000000000000000000000",
2305 => "000000000000000000000000",
2306 => "000000000000000000000000",
2307 => "000000000000000000000000",
2308 => "000000000000000000000000",
2309 => "000000000000000000000000",
2310 => "000000000000000000000000",
2311 => "000000000000000000000000",
2312 => "000000000000000000000000",
2313 => "000000000000000000000000",
2314 => "000000000000000000000000",
2315 => "000000000000000000000000",
2316 => "000000000000000000000000",
2317 => "000000100000001000000010",
2318 => "010000110100001101000011",
2319 => "010000110100001101000011",
2320 => "000101010001010100010101",
2321 => "000000000000000000000000",
2322 => "000000000000000000000000",
2323 => "000000000000000000000000",
2324 => "000000000000000000000000",
2325 => "000000000000000000000000",
2326 => "000000000000000000000000",
2327 => "000000000000000000000000",
2328 => "000000000000000000000000",
2329 => "000000000000000000000000",
2330 => "000000000000000000000000",
2331 => "000000000000000000000000",
2332 => "000000000000000000000000",
2333 => "000000000000000000000000",
2334 => "000000000000000000000000",
2335 => "000000000000000000000000",
2336 => "000000000000000000000000",
2337 => "000000000000000000000000",
2338 => "000000000000000000000000",
2339 => "000000000000000000000000",
2340 => "000000000000000000000000",
2341 => "000000000000000000000000",
2342 => "000000000000000000000000",
2343 => "000000000000000000000000",
2344 => "000000000000000000000000",
2345 => "000000000000000000000000",
2346 => "000000000000000000000000",
2347 => "000000000000000000000000",
2348 => "000000000000000000000000",
2349 => "000000000000000000000000",
2350 => "000000000000000000000000",
2351 => "000000000000000000000000",
2352 => "000000000000000000000000",
2353 => "000000000000000000000000",
2354 => "000000000000000000000000",
2355 => "000000000000000000000000",
2356 => "000000000000000000000000",
2357 => "000000000000000000000000",
2358 => "000000000000000000000000",
2359 => "000000000000000000000000",
2360 => "000000000000000000000000",
2361 => "000000000000000000000000",
2362 => "000000000000000000000000",
2363 => "000000000000000000000000",
2364 => "000000000000000000000000",
2365 => "000000000000000000000000",
2366 => "000000000000000000000000",
2367 => "000000000000000000000000",
2368 => "000000000000000000000000",
2369 => "000000000000000000000000",
2370 => "000000000000000000000000",
2371 => "000000000000000000000000",
2372 => "000000000000000000000000",
2373 => "000000000000000000000000",
2374 => "000000000000000000000000",
2375 => "000000000000000000000000",
2376 => "000000000000000000000000",
2377 => "000000000000000000000000",
2378 => "000000000000000000000000",
2379 => "000000000000000000000000",
2380 => "000000000000000000000000",
2381 => "000000000000000000000000",
2382 => "000000000000000000000000",
2383 => "000000000000000000000000",
2384 => "000000000000000000000000",
2385 => "000000000000000000000000",
2386 => "000000000000000000000000",
2387 => "000000000000000000000000",
2388 => "000000000000000000000000",
2389 => "000000000000000000000000",
2390 => "000000000000000000000000",
2391 => "000000000000000000000000",
2392 => "000000000000000000000000",
2393 => "000000000000000000000000",
2394 => "000000000000000000000000",
2395 => "000000000000000000000000",
2396 => "000000000000000000000000",
2397 => "000000000000000000000000",
2398 => "000000000000000000000000",
2399 => "000000000000000000000000",
2400 => "000000000000000000000000",
2401 => "000000000000000000000000",
2402 => "000000000000000000000000",
2403 => "000000000000000000000000",
2404 => "000000000000000000000000",
2405 => "000000000000000000000000",
2406 => "000000000000000000000000",
2407 => "000000000000000000000000",
2408 => "000000000000000000000000",
2409 => "000000000000000000000000",
2410 => "000000000000000000000000",
2411 => "000000000000000000000000",
2412 => "000000000000000000000000",
2413 => "000000000000000000000000",
2414 => "000000000000000000000000",
2415 => "000000000000000000000000",
2416 => "000000000000000000000000",
2417 => "000000000000000000000000",
2418 => "000000000000000000000000",
2419 => "000000000000000000000000",
2420 => "000000000000000000000000",
2421 => "000000000000000000000000",
2422 => "000000000000000000000000",
2423 => "000000000000000000000000",
2424 => "000000000000000000000000",
2425 => "000000000000000000000000",
2426 => "000000000000000000000000",
2427 => "000000000000000000000000",
2428 => "000000000000000000000000",
2429 => "000000000000000000000000",
2430 => "000000000000000000000000",
2431 => "000000000000000000000000",
2432 => "000000000000000000000000",
2433 => "000000000000000000000000",
2434 => "000000000000000000000000",
2435 => "000000000000000000000000",
2436 => "000000000000000000000000",
2437 => "000000000000000000000000",
2438 => "000000000000000000000000",
2439 => "000000000000000000000000",
2440 => "000000000000000000000000",
2441 => "000000000000000000000000",
2442 => "000000000000000000000000",
2443 => "000000000000000000000000",
2444 => "000000000000000000000000",
2445 => "000000000000000000000000",
2446 => "000000000000000000000000",
2447 => "000000000000000000000000",
2448 => "000000000000000000000000",
2449 => "000000000000000000000000",
2450 => "000000000000000000000000",
2451 => "000000000000000000000000",
2452 => "000000000000000000000000",
2453 => "000000000000000000000000",
2454 => "000000000000000000000000",
2455 => "000000000000000000000000",
2456 => "000000000000000000000000",
2457 => "000000000000000000000000",
2458 => "000000000000000000000000",
2459 => "000000000000000000000000",
2460 => "000000000000000000000000",
2461 => "000000000000000000000000",
2462 => "000000000000000000000000",
2463 => "000000000000000000000000",
2464 => "000000000000000000000000",
2465 => "000000000000000000000000",
2466 => "000000000000000000000000",
2467 => "000000100000001000000010",
2468 => "010000110100001101000011",
2469 => "010000110100001101000011",
2470 => "000101010001010100010101",
2471 => "000000000000000000000000",
2472 => "000000000000000000000000",
2473 => "000000000000000000000000",
2474 => "000000000000000000000000",
2475 => "000000000000000000000000",
2476 => "000000000000000000000000",
2477 => "000000000000000000000000",
2478 => "000000000000000000000000",
2479 => "000000000000000000000000",
2480 => "000000000000000000000000",
2481 => "000000000000000000000000",
2482 => "000000000000000000000000",
2483 => "000000000000000000000000",
2484 => "000000000000000000000000",
2485 => "000000000000000000000000",
2486 => "000000000000000000000000",
2487 => "000000000000000000000000",
2488 => "000000000000000000000000",
2489 => "000000000000000000000000",
2490 => "000000000000000000000000",
2491 => "000000000000000000000000",
2492 => "000000000000000000000000",
2493 => "000000000000000000000000",
2494 => "000000000000000000000000",
2495 => "000000000000000000000000",
2496 => "000000000000000000000000",
2497 => "000000000000000000000000",
2498 => "000000000000000000000000",
2499 => "000000000000000000000000",
2500 => "000000000000000000000000",
2501 => "000000000000000000000000",
2502 => "000000000000000000000000",
2503 => "000000000000000000000000",
2504 => "000000000000000000000000",
2505 => "000000000000000000000000",
2506 => "000000000000000000000000",
2507 => "000000000000000000000000",
2508 => "000000000000000000000000",
2509 => "000000000000000000000000",
2510 => "000000000000000000000000",
2511 => "000000000000000000000000",
2512 => "000000000000000000000000",
2513 => "000000000000000000000000",
2514 => "000000000000000000000000",
2515 => "000000000000000000000000",
2516 => "000000000000000000000000",
2517 => "000000000000000000000000",
2518 => "000000000000000000000000",
2519 => "000000000000000000000000",
2520 => "000000000000000000000000",
2521 => "000000000000000000000000",
2522 => "000000000000000000000000",
2523 => "000000000000000000000000",
2524 => "000000000000000000000000",
2525 => "000000000000000000000000",
2526 => "000000000000000000000000",
2527 => "000000000000000000000000",
2528 => "000000000000000000000000",
2529 => "000000000000000000000000",
2530 => "000000000000000000000000",
2531 => "000000000000000000000000",
2532 => "000000000000000000000000",
2533 => "000000000000000000000000",
2534 => "000000000000000000000000",
2535 => "000000000000000000000000",
2536 => "000000000000000000000000",
2537 => "000000000000000000000000",
2538 => "000000000000000000000000",
2539 => "000000000000000000000000",
2540 => "000000000000000000000000",
2541 => "000000000000000000000000",
2542 => "000000000000000000000000",
2543 => "000000000000000000000000",
2544 => "000000000000000000000000",
2545 => "000000000000000000000000",
2546 => "000000000000000000000000",
2547 => "000000000000000000000000",
2548 => "000000000000000000000000",
2549 => "000000000000000000000000",
2550 => "000000000000000000000000",
2551 => "000000000000000000000000",
2552 => "000000000000000000000000",
2553 => "000000000000000000000000",
2554 => "000000000000000000000000",
2555 => "000000000000000000000000",
2556 => "000000000000000000000000",
2557 => "000000000000000000000000",
2558 => "000000000000000000000000",
2559 => "000000000000000000000000",
2560 => "000000000000000000000000",
2561 => "000000000000000000000000",
2562 => "000000000000000000000000",
2563 => "000000000000000000000000",
2564 => "000000000000000000000000",
2565 => "000000000000000000000000",
2566 => "000000000000000000000000",
2567 => "000000000000000000000000",
2568 => "000000000000000000000000",
2569 => "000000000000000000000000",
2570 => "000000000000000000000000",
2571 => "000000000000000000000000",
2572 => "000000000000000000000000",
2573 => "000000000000000000000000",
2574 => "000000000000000000000000",
2575 => "000000000000000000000000",
2576 => "000000000000000000000000",
2577 => "000000000000000000000000",
2578 => "000000000000000000000000",
2579 => "000000000000000000000000",
2580 => "000000000000000000000000",
2581 => "000000000000000000000000",
2582 => "000000000000000000000000",
2583 => "000000000000000000000000",
2584 => "000000000000000000000000",
2585 => "000000000000000000000000",
2586 => "000000000000000000000000",
2587 => "000000000000000000000000",
2588 => "000000000000000000000000",
2589 => "000000000000000000000000",
2590 => "000000000000000000000000",
2591 => "000000000000000000000000",
2592 => "000000000000000000000000",
2593 => "000000000000000000000000",
2594 => "000000000000000000000000",
2595 => "000000000000000000000000",
2596 => "000000000000000000000000",
2597 => "000000000000000000000000",
2598 => "000000000000000000000000",
2599 => "000000000000000000000000",
2600 => "000000000000000000000000",
2601 => "000000000000000000000000",
2602 => "000000000000000000000000",
2603 => "000000000000000000000000",
2604 => "000000000000000000000000",
2605 => "000000000000000000000000",
2606 => "000000000000000000000000",
2607 => "000000000000000000000000",
2608 => "000000000000000000000000",
2609 => "000000000000000000000000",
2610 => "000000000000000000000000",
2611 => "000000000000000000000000",
2612 => "000000000000000000000000",
2613 => "000000000000000000000000",
2614 => "000000000000000000000000",
2615 => "000000000000000000000000",
2616 => "000000000000000000000000",
2617 => "000000100000001000000010",
2618 => "010000110100001101000011",
2619 => "010000110100001101000011",
2620 => "000101010001010100010101",
2621 => "000000000000000000000000",
2622 => "000000000000000000000000",
2623 => "000000000000000000000000",
2624 => "000000000000000000000000",
2625 => "000000000000000000000000",
2626 => "000000000000000000000000",
2627 => "000000000000000000000000",
2628 => "000000000000000000000000",
2629 => "000000000000000000000000",
2630 => "000000000000000000000000",
2631 => "000000000000000000000000",
2632 => "000000000000000000000000",
2633 => "000000000000000000000000",
2634 => "000000000000000000000000",
2635 => "000000000000000000000000",
2636 => "000000000000000000000000",
2637 => "000000000000000000000000",
2638 => "000000000000000000000000",
2639 => "000000000000000000000000",
2640 => "000000000000000000000000",
2641 => "000000000000000000000000",
2642 => "000000000000000000000000",
2643 => "000000000000000000000000",
2644 => "000000000000000000000000",
2645 => "000000000000000000000000",
2646 => "000000000000000000000000",
2647 => "000000000000000000000000",
2648 => "000000000000000000000000",
2649 => "000000000000000000000000",
2650 => "000000000000000000000000",
2651 => "000000000000000000000000",
2652 => "000000000000000000000000",
2653 => "000000000000000000000000",
2654 => "000000000000000000000000",
2655 => "000000000000000000000000",
2656 => "000000000000000000000000",
2657 => "000000000000000000000000",
2658 => "000000000000000000000000",
2659 => "000000000000000000000000",
2660 => "000000000000000000000000",
2661 => "000000000000000000000000",
2662 => "000000000000000000000000",
2663 => "000000000000000000000000",
2664 => "000000000000000000000000",
2665 => "000000000000000000000000",
2666 => "000000000000000000000000",
2667 => "000000000000000000000000",
2668 => "000000000000000000000000",
2669 => "000000000000000000000000",
2670 => "000000000000000000000000",
2671 => "000000000000000000000000",
2672 => "000000000000000000000000",
2673 => "000000000000000000000000",
2674 => "000000000000000000000000",
2675 => "000000000000000000000000",
2676 => "000000000000000000000000",
2677 => "000000000000000000000000",
2678 => "000000000000000000000000",
2679 => "000000000000000000000000",
2680 => "000000000000000000000000",
2681 => "000000000000000000000000",
2682 => "000000000000000000000000",
2683 => "000000000000000000000000",
2684 => "000000000000000000000000",
2685 => "000000000000000000000000",
2686 => "000000000000000000000000",
2687 => "000000000000000000000000",
2688 => "000000000000000000000000",
2689 => "000000000000000000000000",
2690 => "000000000000000000000000",
2691 => "000000000000000000000000",
2692 => "000000000000000000000000",
2693 => "000000000000000000000000",
2694 => "000000000000000000000000",
2695 => "000000000000000000000000",
2696 => "000000000000000000000000",
2697 => "000000000000000000000000",
2698 => "000000000000000000000000",
2699 => "000000000000000000000000",
2700 => "000000000000000000000000",
2701 => "000000000000000000000000",
2702 => "000000000000000000000000",
2703 => "000000000000000000000000",
2704 => "000000000000000000000000",
2705 => "000000000000000000000000",
2706 => "000000000000000000000000",
2707 => "000000000000000000000000",
2708 => "000000000000000000000000",
2709 => "000000000000000000000000",
2710 => "000000000000000000000000",
2711 => "000000000000000000000000",
2712 => "000000000000000000000000",
2713 => "000000000000000000000000",
2714 => "000000000000000000000000",
2715 => "000000000000000000000000",
2716 => "000000000000000000000000",
2717 => "000000000000000000000000",
2718 => "000000000000000000000000",
2719 => "000000000000000000000000",
2720 => "000000000000000000000000",
2721 => "000000000000000000000000",
2722 => "000000000000000000000000",
2723 => "000000000000000000000000",
2724 => "000000000000000000000000",
2725 => "000000000000000000000000",
2726 => "000000000000000000000000",
2727 => "000000000000000000000000",
2728 => "000000000000000000000000",
2729 => "000000000000000000000000",
2730 => "000000000000000000000000",
2731 => "000000000000000000000000",
2732 => "000000000000000000000000",
2733 => "000000000000000000000000",
2734 => "000000000000000000000000",
2735 => "000000000000000000000000",
2736 => "000000000000000000000000",
2737 => "000000000000000000000000",
2738 => "000000000000000000000000",
2739 => "000000000000000000000000",
2740 => "000000000000000000000000",
2741 => "000000000000000000000000",
2742 => "000000000000000000000000",
2743 => "000000000000000000000000",
2744 => "000000000000000000000000",
2745 => "000000000000000000000000",
2746 => "000000000000000000000000",
2747 => "000000000000000000000000",
2748 => "000000000000000000000000",
2749 => "000000000000000000000000",
2750 => "000000000000000000000000",
2751 => "000000000000000000000000",
2752 => "000000000000000000000000",
2753 => "000000000000000000000000",
2754 => "000000000000000000000000",
2755 => "000000000000000000000000",
2756 => "000000000000000000000000",
2757 => "000000000000000000000000",
2758 => "000000000000000000000000",
2759 => "000000000000000000000000",
2760 => "000000000000000000000000",
2761 => "000000000000000000000000",
2762 => "000000000000000000000000",
2763 => "000000000000000000000000",
2764 => "000000000000000000000000",
2765 => "000001100000011000000110",
2766 => "000100010001000100010001",
2767 => "000100100001001000010010",
2768 => "010000110100001101000011",
2769 => "010000110100001101000011",
2770 => "001000000010000000100000",
2771 => "000100010001000100010001",
2772 => "000010110000101100001011",
2773 => "000000000000000000000000",
2774 => "000000000000000000000000",
2775 => "000000000000000000000000",
2776 => "000000000000000000000000",
2777 => "000000000000000000000000",
2778 => "000000000000000000000000",
2779 => "000000000000000000000000",
2780 => "000000000000000000000000",
2781 => "000000000000000000000000",
2782 => "000000000000000000000000",
2783 => "000000000000000000000000",
2784 => "000000000000000000000000",
2785 => "000000000000000000000000",
2786 => "000000000000000000000000",
2787 => "000000000000000000000000",
2788 => "000000000000000000000000",
2789 => "000000000000000000000000",
2790 => "000000000000000000000000",
2791 => "000000000000000000000000",
2792 => "000000000000000000000000",
2793 => "000000000000000000000000",
2794 => "000000000000000000000000",
2795 => "000000000000000000000000",
2796 => "000000000000000000000000",
2797 => "000000000000000000000000",
2798 => "000000000000000000000000",
2799 => "000000000000000000000000",
2800 => "000000000000000000000000",
2801 => "000000000000000000000000",
2802 => "000000000000000000000000",
2803 => "000000000000000000000000",
2804 => "000000000000000000000000",
2805 => "000000000000000000000000",
2806 => "000000000000000000000000",
2807 => "000000000000000000000000",
2808 => "000000000000000000000000",
2809 => "000000000000000000000000",
2810 => "000000000000000000000000",
2811 => "000000000000000000000000",
2812 => "000000000000000000000000",
2813 => "000000000000000000000000",
2814 => "000000000000000000000000",
2815 => "000000000000000000000000",
2816 => "000000000000000000000000",
2817 => "000000000000000000000000",
2818 => "000000000000000000000000",
2819 => "000000000000000000000000",
2820 => "000000000000000000000000",
2821 => "000000000000000000000000",
2822 => "000000000000000000000000",
2823 => "000000000000000000000000",
2824 => "000000000000000000000000",
2825 => "000000000000000000000000",
2826 => "000000000000000000000000",
2827 => "000000000000000000000000",
2828 => "000000000000000000000000",
2829 => "000000000000000000000000",
2830 => "000000000000000000000000",
2831 => "000000000000000000000000",
2832 => "000000000000000000000000",
2833 => "000000000000000000000000",
2834 => "000000000000000000000000",
2835 => "000000000000000000000000",
2836 => "000000000000000000000000",
2837 => "000000000000000000000000",
2838 => "000000000000000000000000",
2839 => "000000000000000000000000",
2840 => "000000000000000000000000",
2841 => "000000000000000000000000",
2842 => "000000000000000000000000",
2843 => "000000000000000000000000",
2844 => "000000000000000000000000",
2845 => "000000000000000000000000",
2846 => "000000000000000000000000",
2847 => "000000000000000000000000",
2848 => "000000000000000000000000",
2849 => "000000000000000000000000",
2850 => "000000000000000000000000",
2851 => "000000000000000000000000",
2852 => "000000000000000000000000",
2853 => "000000000000000000000000",
2854 => "000000000000000000000000",
2855 => "000000000000000000000000",
2856 => "000000000000000000000000",
2857 => "000000000000000000000000",
2858 => "000000000000000000000000",
2859 => "000000000000000000000000",
2860 => "000000000000000000000000",
2861 => "000000000000000000000000",
2862 => "000000000000000000000000",
2863 => "000000000000000000000000",
2864 => "000000000000000000000000",
2865 => "000000000000000000000000",
2866 => "000000000000000000000000",
2867 => "000000000000000000000000",
2868 => "000000000000000000000000",
2869 => "000000000000000000000000",
2870 => "000000000000000000000000",
2871 => "000000000000000000000000",
2872 => "000000000000000000000000",
2873 => "000000000000000000000000",
2874 => "000000000000000000000000",
2875 => "000000000000000000000000",
2876 => "000000000000000000000000",
2877 => "000000000000000000000000",
2878 => "000000000000000000000000",
2879 => "000000000000000000000000",
2880 => "000000000000000000000000",
2881 => "000000000000000000000000",
2882 => "000000000000000000000000",
2883 => "000000000000000000000000",
2884 => "000000000000000000000000",
2885 => "000000000000000000000000",
2886 => "000000000000000000000000",
2887 => "000000000000000000000000",
2888 => "000000000000000000000000",
2889 => "000000000000000000000000",
2890 => "000000000000000000000000",
2891 => "000000000000000000000000",
2892 => "000000000000000000000000",
2893 => "000000000000000000000000",
2894 => "000000000000000000000000",
2895 => "000000000000000000000000",
2896 => "000000000000000000000000",
2897 => "000000000000000000000000",
2898 => "000000000000000000000000",
2899 => "000000000000000000000000",
2900 => "000000000000000000000000",
2901 => "000000000000000000000000",
2902 => "000000000000000000000000",
2903 => "000000000000000000000000",
2904 => "000000000000000000000000",
2905 => "000000000000000000000000",
2906 => "000000000000000000000000",
2907 => "000000000000000000000000",
2908 => "000000000000000000000000",
2909 => "000000000000000000000000",
2910 => "000000000000000000000000",
2911 => "000000000000000000000000",
2912 => "000000000000000000000000",
2913 => "000000000000000000000000",
2914 => "000000000000000000000000",
2915 => "000110010001100100011001",
2916 => "010000110100001101000011",
2917 => "010000110100001101000011",
2918 => "010000110100001101000011",
2919 => "010000110100001101000011",
2920 => "010000110100001101000011",
2921 => "010000110100001101000011",
2922 => "001011000010110000101100",
2923 => "000000000000000000000000",
2924 => "000000000000000000000000",
2925 => "000000000000000000000000",
2926 => "000000000000000000000000",
2927 => "000000000000000000000000",
2928 => "000000000000000000000000",
2929 => "000000000000000000000000",
2930 => "000000000000000000000000",
2931 => "000000000000000000000000",
2932 => "000000000000000000000000",
2933 => "000000000000000000000000",
2934 => "000000000000000000000000",
2935 => "000000000000000000000000",
2936 => "000000000000000000000000",
2937 => "000000000000000000000000",
2938 => "000000000000000000000000",
2939 => "000000000000000000000000",
2940 => "000000000000000000000000",
2941 => "000000000000000000000000",
2942 => "000000000000000000000000",
2943 => "000000000000000000000000",
2944 => "000000000000000000000000",
2945 => "000000000000000000000000",
2946 => "000000000000000000000000",
2947 => "000000000000000000000000",
2948 => "000000000000000000000000",
2949 => "000000000000000000000000",
2950 => "000000000000000000000000",
2951 => "000000000000000000000000",
2952 => "000000000000000000000000",
2953 => "000000000000000000000000",
2954 => "000000000000000000000000",
2955 => "000000000000000000000000",
2956 => "000000000000000000000000",
2957 => "000000000000000000000000",
2958 => "000000000000000000000000",
2959 => "000000000000000000000000",
2960 => "000000000000000000000000",
2961 => "000000000000000000000000",
2962 => "000000000000000000000000",
2963 => "000000000000000000000000",
2964 => "000000000000000000000000",
2965 => "000000000000000000000000",
2966 => "000000000000000000000000",
2967 => "000000000000000000000000",
2968 => "000000000000000000000000",
2969 => "000000000000000000000000",
2970 => "000000000000000000000000",
2971 => "000000000000000000000000",
2972 => "000000000000000000000000",
2973 => "000000000000000000000000",
2974 => "000000000000000000000000",
2975 => "000000000000000000000000",
2976 => "000000000000000000000000",
2977 => "000000000000000000000000",
2978 => "000000000000000000000000",
2979 => "000000000000000000000000",
2980 => "000000000000000000000000",
2981 => "000000000000000000000000",
2982 => "000000000000000000000000",
2983 => "000000000000000000000000",
2984 => "000000000000000000000000",
2985 => "000000000000000000000000",
2986 => "000000000000000000000000",
2987 => "000000000000000000000000",
2988 => "000000000000000000000000",
2989 => "000000000000000000000000",
2990 => "000000000000000000000000",
2991 => "000000000000000000000000",
2992 => "000000000000000000000000",
2993 => "000000000000000000000000",
2994 => "000000000000000000000000",
2995 => "000000000000000000000000",
2996 => "000000000000000000000000",
2997 => "000000000000000000000000",
2998 => "000000000000000000000000",
2999 => "000000000000000000000000",
3000 => "000000000000000000000000",
3001 => "000000000000000000000000",
3002 => "000000000000000000000000",
3003 => "000000000000000000000000",
3004 => "000000000000000000000000",
3005 => "000000000000000000000000",
3006 => "000000000000000000000000",
3007 => "000000000000000000000000",
3008 => "000000000000000000000000",
3009 => "000000000000000000000000",
3010 => "000000000000000000000000",
3011 => "000000000000000000000000",
3012 => "000000000000000000000000",
3013 => "000000000000000000000000",
3014 => "000000000000000000000000",
3015 => "000000000000000000000000",
3016 => "000000000000000000000000",
3017 => "000000000000000000000000",
3018 => "000000000000000000000000",
3019 => "000000000000000000000000",
3020 => "000000000000000000000000",
3021 => "000000000000000000000000",
3022 => "000000000000000000000000",
3023 => "000000000000000000000000",
3024 => "000000000000000000000000",
3025 => "000000000000000000000000",
3026 => "000000000000000000000000",
3027 => "000000000000000000000000",
3028 => "000000000000000000000000",
3029 => "000000000000000000000000",
3030 => "000000000000000000000000",
3031 => "000000000000000000000000",
3032 => "000000000000000000000000",
3033 => "000000000000000000000000",
3034 => "000000000000000000000000",
3035 => "000000000000000000000000",
3036 => "000000000000000000000000",
3037 => "000000000000000000000000",
3038 => "000000000000000000000000",
3039 => "000000000000000000000000",
3040 => "000000000000000000000000",
3041 => "000000000000000000000000",
3042 => "000000000000000000000000",
3043 => "000000000000000000000000",
3044 => "000000000000000000000000",
3045 => "000000000000000000000000",
3046 => "000000000000000000000000",
3047 => "000000000000000000000000",
3048 => "000000000000000000000000",
3049 => "000000000000000000000000",
3050 => "000000000000000000000000",
3051 => "000000000000000000000000",
3052 => "000000000000000000000000",
3053 => "000000000000000000000000",
3054 => "000000000000000000000000",
3055 => "000000000000000000000000",
3056 => "000000000000000000000000",
3057 => "000000000000000000000000",
3058 => "000000000000000000000000",
3059 => "000000000000000000000000",
3060 => "000000000000000000000000",
3061 => "000000000000000000000000",
3062 => "000000000000000000000000",
3063 => "000000000000000000000000",
3064 => "000000000000000000000000",
3065 => "000110010001100100011001",
3066 => "010000110100001101000011",
3067 => "010000110100001101000011",
3068 => "010000110100001101000011",
3069 => "010000110100001101000011",
3070 => "010000110100001101000011",
3071 => "010000110100001101000011",
3072 => "001011000010110000101100",
3073 => "000000000000000000000000",
3074 => "000000000000000000000000",
3075 => "000000000000000000000000",
3076 => "000000000000000000000000",
3077 => "000000000000000000000000",
3078 => "000000000000000000000000",
3079 => "000000000000000000000000",
3080 => "000000000000000000000000",
3081 => "000000000000000000000000",
3082 => "000000000000000000000000",
3083 => "000000000000000000000000",
3084 => "000000000000000000000000",
3085 => "000000000000000000000000",
3086 => "000000000000000000000000",
3087 => "000000000000000000000000",
3088 => "000000000000000000000000",
3089 => "000000000000000000000000",
3090 => "000000000000000000000000",
3091 => "000000000000000000000000",
3092 => "000000000000000000000000",
3093 => "000000000000000000000000",
3094 => "000000000000000000000000",
3095 => "000000000000000000000000",
3096 => "000000000000000000000000",
3097 => "000000000000000000000000",
3098 => "000000000000000000000000",
3099 => "000000000000000000000000",
3100 => "000000000000000000000000",
3101 => "000000000000000000000000",
3102 => "000000000000000000000000",
3103 => "000000000000000000000000",
3104 => "000000000000000000000000",
3105 => "000000000000000000000000",
3106 => "000000000000000000000000",
3107 => "000000000000000000000000",
3108 => "000000000000000000000000",
3109 => "000000000000000000000000",
3110 => "000000000000000000000000",
3111 => "000000000000000000000000",
3112 => "000000000000000000000000",
3113 => "000000000000000000000000",
3114 => "000000000000000000000000",
3115 => "000000000000000000000000",
3116 => "000000000000000000000000",
3117 => "000000000000000000000000",
3118 => "000000000000000000000000",
3119 => "000000000000000000000000",
3120 => "000000000000000000000000",
3121 => "000000000000000000000000",
3122 => "000000000000000000000000",
3123 => "000000000000000000000000",
3124 => "000000000000000000000000",
3125 => "000000000000000000000000",
3126 => "000000000000000000000000",
3127 => "000000000000000000000000",
3128 => "000000000000000000000000",
3129 => "000000000000000000000000",
3130 => "000000000000000000000000",
3131 => "000000000000000000000000",
3132 => "000000000000000000000000",
3133 => "000000000000000000000000",
3134 => "000000000000000000000000",
3135 => "000000000000000000000000",
3136 => "000000000000000000000000",
3137 => "000000000000000000000000",
3138 => "000000000000000000000000",
3139 => "000000000000000000000000",
3140 => "000000000000000000000000",
3141 => "000000000000000000000000",
3142 => "000000000000000000000000",
3143 => "000000000000000000000000",
3144 => "000000000000000000000000",
3145 => "000000000000000000000000",
3146 => "000000000000000000000000",
3147 => "000000000000000000000000",
3148 => "000000000000000000000000",
3149 => "000000000000000000000000",
3150 => "000000000000000000000000",
3151 => "000000000000000000000000",
3152 => "000000000000000000000000",
3153 => "000000000000000000000000",
3154 => "000000000000000000000000",
3155 => "000000000000000000000000",
3156 => "000000000000000000000000",
3157 => "000000000000000000000000",
3158 => "000000000000000000000000",
3159 => "000000000000000000000000",
3160 => "000000000000000000000000",
3161 => "000000000000000000000000",
3162 => "000000000000000000000000",
3163 => "000000000000000000000000",
3164 => "000000000000000000000000",
3165 => "000000000000000000000000",
3166 => "000000000000000000000000",
3167 => "000000000000000000000000",
3168 => "000000000000000000000000",
3169 => "000000000000000000000000",
3170 => "000000000000000000000000",
3171 => "000000000000000000000000",
3172 => "000000000000000000000000",
3173 => "000000000000000000000000",
3174 => "000000000000000000000000",
3175 => "000000000000000000000000",
3176 => "000000000000000000000000",
3177 => "000000000000000000000000",
3178 => "000000000000000000000000",
3179 => "000000000000000000000000",
3180 => "000000000000000000000000",
3181 => "000000000000000000000000",
3182 => "000000000000000000000000",
3183 => "000000000000000000000000",
3184 => "000000000000000000000000",
3185 => "000000000000000000000000",
3186 => "000000000000000000000000",
3187 => "000000000000000000000000",
3188 => "000000000000000000000000",
3189 => "000000000000000000000000",
3190 => "000000000000000000000000",
3191 => "000000000000000000000000",
3192 => "000000000000000000000000",
3193 => "000000000000000000000000",
3194 => "000000000000000000000000",
3195 => "000000000000000000000000",
3196 => "000000000000000000000000",
3197 => "000000000000000000000000",
3198 => "000000000000000000000000",
3199 => "000000000000000000000000",
3200 => "000000000000000000000000",
3201 => "000000000000000000000000",
3202 => "000000000000000000000000",
3203 => "000000000000000000000000",
3204 => "000000000000000000000000",
3205 => "000000000000000000000000",
3206 => "000000000000000000000000",
3207 => "000000000000000000000000",
3208 => "000000000000000000000000",
3209 => "000000000000000000000000",
3210 => "000000000000000000000000",
3211 => "000000000000000000000000",
3212 => "000000000000000000000000",
3213 => "000000000000000000000000",
3214 => "000000000000000000000000",
3215 => "000110010001100100011001",
3216 => "010000110100001101000011",
3217 => "010000110100001101000011",
3218 => "010000110100001101000011",
3219 => "010000110100001101000011",
3220 => "010000110100001101000011",
3221 => "010000110100001101000011",
3222 => "001011000010110000101100",
3223 => "000000000000000000000000",
3224 => "000000000000000000000000",
3225 => "000000000000000000000000",
3226 => "000000000000000000000000",
3227 => "000000000000000000000000",
3228 => "000000000000000000000000",
3229 => "000000000000000000000000",
3230 => "000000000000000000000000",
3231 => "000000000000000000000000",
3232 => "000000000000000000000000",
3233 => "000000000000000000000000",
3234 => "000000000000000000000000",
3235 => "000000000000000000000000",
3236 => "000000000000000000000000",
3237 => "000000000000000000000000",
3238 => "000000000000000000000000",
3239 => "000000000000000000000000",
3240 => "000000000000000000000000",
3241 => "000000000000000000000000",
3242 => "000000000000000000000000",
3243 => "000000000000000000000000",
3244 => "000000000000000000000000",
3245 => "000000000000000000000000",
3246 => "000000000000000000000000",
3247 => "000000000000000000000000",
3248 => "000000000000000000000000",
3249 => "000000000000000000000000",
3250 => "000000000000000000000000",
3251 => "000000000000000000000000",
3252 => "000000000000000000000000",
3253 => "000000000000000000000000",
3254 => "000000000000000000000000",
3255 => "000000000000000000000000",
3256 => "000000000000000000000000",
3257 => "000000000000000000000000",
3258 => "000000000000000000000000",
3259 => "000000000000000000000000",
3260 => "000000000000000000000000",
3261 => "000000000000000000000000",
3262 => "000000000000000000000000",
3263 => "000000000000000000000000",
3264 => "000000000000000000000000",
3265 => "000000000000000000000000",
3266 => "000000000000000000000000",
3267 => "000000000000000000000000",
3268 => "000000000000000000000000",
3269 => "000000000000000000000000",
3270 => "000000000000000000000000",
3271 => "000000000000000000000000",
3272 => "000000000000000000000000",
3273 => "000000000000000000000000",
3274 => "000000000000000000000000",
3275 => "000000000000000000000000",
3276 => "000000000000000000000000",
3277 => "000000000000000000000000",
3278 => "000000000000000000000000",
3279 => "000000000000000000000000",
3280 => "000000000000000000000000",
3281 => "000000000000000000000000",
3282 => "000000000000000000000000",
3283 => "000000000000000000000000",
3284 => "000000000000000000000000",
3285 => "000000000000000000000000",
3286 => "000000000000000000000000",
3287 => "000000000000000000000000",
3288 => "000000000000000000000000",
3289 => "000000000000000000000000",
3290 => "000000000000000000000000",
3291 => "000000000000000000000000",
3292 => "000000000000000000000000",
3293 => "000000000000000000000000",
3294 => "000000000000000000000000",
3295 => "000000000000000000000000",
3296 => "000000000000000000000000",
3297 => "000000000000000000000000",
3298 => "000000000000000000000000",
3299 => "000000000000000000000000",
3300 => "000000000000000000000000",
3301 => "000000000000000000000000",
3302 => "000000000000000000000000",
3303 => "000000000000000000000000",
3304 => "000000000000000000000000",
3305 => "000000000000000000000000",
3306 => "000000000000000000000000",
3307 => "000000000000000000000000",
3308 => "000000000000000000000000",
3309 => "000000000000000000000000",
3310 => "000000000000000000000000",
3311 => "000000000000000000000000",
3312 => "000000000000000000000000",
3313 => "000000000000000000000000",
3314 => "000000000000000000000000",
3315 => "000000000000000000000000",
3316 => "000000000000000000000000",
3317 => "000000000000000000000000",
3318 => "000000000000000000000000",
3319 => "000000000000000000000000",
3320 => "000000000000000000000000",
3321 => "000000000000000000000000",
3322 => "000000000000000000000000",
3323 => "000000000000000000000000",
3324 => "000000000000000000000000",
3325 => "000000000000000000000000",
3326 => "000000000000000000000000",
3327 => "000000000000000000000000",
3328 => "000000000000000000000000",
3329 => "000000000000000000000000",
3330 => "000000000000000000000000",
3331 => "000000000000000000000000",
3332 => "000000000000000000000000",
3333 => "000000000000000000000000",
3334 => "000000000000000000000000",
3335 => "000000000000000000000000",
3336 => "000000000000000000000000",
3337 => "000000000000000000000000",
3338 => "000000000000000000000000",
3339 => "000000000000000000000000",
3340 => "000000000000000000000000",
3341 => "000000000000000000000000",
3342 => "000000000000000000000000",
3343 => "000000000000000000000000",
3344 => "000000000000000000000000",
3345 => "000000000000000000000000",
3346 => "000000000000000000000000",
3347 => "000000000000000000000000",
3348 => "000000000000000000000000",
3349 => "000000000000000000000000",
3350 => "000000000000000000000000",
3351 => "000000000000000000000000",
3352 => "000000000000000000000000",
3353 => "000000000000000000000000",
3354 => "000000000000000000000000",
3355 => "000000000000000000000000",
3356 => "000000000000000000000000",
3357 => "000000000000000000000000",
3358 => "000000000000000000000000",
3359 => "000000000000000000000000",
3360 => "000000000000000000000000",
3361 => "000000000000000000000000",
3362 => "000000000000000000000000",
3363 => "000000000000000000000000",
3364 => "000000000000000000000000",
3365 => "000110010001100100011001",
3366 => "010000110100001101000011",
3367 => "010000110100001101000011",
3368 => "010000110100001101000011",
3369 => "010000110100001101000011",
3370 => "010000110100001101000011",
3371 => "010000110100001101000011",
3372 => "001011000010110000101100",
3373 => "000000000000000000000000",
3374 => "000000000000000000000000",
3375 => "000000000000000000000000",
3376 => "000000000000000000000000",
3377 => "000000000000000000000000",
3378 => "000000000000000000000000",
3379 => "000000000000000000000000",
3380 => "000000000000000000000000",
3381 => "000000000000000000000000",
3382 => "000000000000000000000000",
3383 => "000000000000000000000000",
3384 => "000000000000000000000000",
3385 => "000000000000000000000000",
3386 => "000000000000000000000000",
3387 => "000000000000000000000000",
3388 => "000000000000000000000000",
3389 => "000000000000000000000000",
3390 => "000000000000000000000000",
3391 => "000000000000000000000000",
3392 => "000000000000000000000000",
3393 => "000000000000000000000000",
3394 => "000000000000000000000000",
3395 => "000000000000000000000000",
3396 => "000000000000000000000000",
3397 => "000000000000000000000000",
3398 => "000000000000000000000000",
3399 => "000000000000000000000000",
3400 => "000000000000000000000000",
3401 => "000000000000000000000000",
3402 => "000000000000000000000000",
3403 => "000000000000000000000000",
3404 => "000000000000000000000000",
3405 => "000000000000000000000000",
3406 => "000000000000000000000000",
3407 => "000000000000000000000000",
3408 => "000000000000000000000000",
3409 => "000000000000000000000000",
3410 => "000000000000000000000000",
3411 => "000000000000000000000000",
3412 => "000000000000000000000000",
3413 => "000000000000000000000000",
3414 => "000000000000000000000000",
3415 => "000000000000000000000000",
3416 => "000000000000000000000000",
3417 => "000000000000000000000000",
3418 => "000000000000000000000000",
3419 => "000000000000000000000000",
3420 => "000000000000000000000000",
3421 => "000000000000000000000000",
3422 => "000000000000000000000000",
3423 => "000000000000000000000000",
3424 => "000000000000000000000000",
3425 => "000000000000000000000000",
3426 => "000000000000000000000000",
3427 => "000000000000000000000000",
3428 => "000000000000000000000000",
3429 => "000000000000000000000000",
3430 => "000000000000000000000000",
3431 => "000000000000000000000000",
3432 => "000000000000000000000000",
3433 => "000000000000000000000000",
3434 => "000000000000000000000000",
3435 => "000000000000000000000000",
3436 => "000000000000000000000000",
3437 => "000000000000000000000000",
3438 => "000000000000000000000000",
3439 => "000000000000000000000000",
3440 => "000000000000000000000000",
3441 => "000000000000000000000000",
3442 => "000000000000000000000000",
3443 => "000000000000000000000000",
3444 => "000000000000000000000000",
3445 => "000000000000000000000000",
3446 => "000000000000000000000000",
3447 => "000000000000000000000000",
3448 => "000000000000000000000000",
3449 => "000000000000000000000000",
3450 => "000000000000000000000000",
3451 => "000000000000000000000000",
3452 => "000000000000000000000000",
3453 => "000000000000000000000000",
3454 => "000000000000000000000000",
3455 => "000000000000000000000000",
3456 => "000000000000000000000000",
3457 => "000000000000000000000000",
3458 => "000000000000000000000000",
3459 => "000000000000000000000000",
3460 => "000000000000000000000000",
3461 => "000000000000000000000000",
3462 => "000000000000000000000000",
3463 => "000000000000000000000000",
3464 => "000000000000000000000000",
3465 => "000000000000000000000000",
3466 => "000000000000000000000000",
3467 => "000000000000000000000000",
3468 => "000000000000000000000000",
3469 => "000000000000000000000000",
3470 => "000000000000000000000000",
3471 => "000000000000000000000000",
3472 => "000000000000000000000000",
3473 => "000000000000000000000000",
3474 => "000000000000000000000000",
3475 => "000000000000000000000000",
3476 => "000000000000000000000000",
3477 => "000000000000000000000000",
3478 => "000000000000000000000000",
3479 => "000000000000000000000000",
3480 => "000000000000000000000000",
3481 => "000000000000000000000000",
3482 => "000000000000000000000000",
3483 => "000000000000000000000000",
3484 => "000000000000000000000000",
3485 => "000000000000000000000000",
3486 => "000000000000000000000000",
3487 => "000000000000000000000000",
3488 => "000000000000000000000000",
3489 => "000000000000000000000000",
3490 => "000000000000000000000000",
3491 => "000000000000000000000000",
3492 => "000000000000000000000000",
3493 => "000000000000000000000000",
3494 => "000000000000000000000000",
3495 => "000000000000000000000000",
3496 => "000000000000000000000000",
3497 => "000000000000000000000000",
3498 => "000000000000000000000000",
3499 => "000000000000000000000000",
3500 => "000000000000000000000000",
3501 => "000000000000000000000000",
3502 => "000000000000000000000000",
3503 => "000000000000000000000000",
3504 => "000000000000000000000000",
3505 => "000000000000000000000000",
3506 => "000000000000000000000000",
3507 => "000000000000000000000000",
3508 => "000000000000000000000000",
3509 => "000000000000000000000000",
3510 => "000000000000000000000000",
3511 => "000000000000000000000000",
3512 => "000000000000000000000000",
3513 => "000000000000000000000000",
3514 => "000000000000000000000000",
3515 => "000110010001100100011001",
3516 => "010000110100001101000011",
3517 => "010000110100001101000011",
3518 => "010000110100001101000011",
3519 => "010000110100001101000011",
3520 => "010000110100001101000011",
3521 => "010000110100001101000011",
3522 => "001011000010110000101100",
3523 => "000000000000000000000000",
3524 => "000000000000000000000000",
3525 => "000000000000000000000000",
3526 => "000000000000000000000000",
3527 => "000000000000000000000000",
3528 => "000000000000000000000000",
3529 => "000000000000000000000000",
3530 => "000000000000000000000000",
3531 => "000000000000000000000000",
3532 => "000000000000000000000000",
3533 => "000000000000000000000000",
3534 => "000000000000000000000000",
3535 => "000000000000000000000000",
3536 => "000000000000000000000000",
3537 => "000000000000000000000000",
3538 => "000000000000000000000000",
3539 => "000000000000000000000000",
3540 => "000000000000000000000000",
3541 => "000000000000000000000000",
3542 => "000000000000000000000000",
3543 => "000000000000000000000000",
3544 => "000000000000000000000000",
3545 => "000000000000000000000000",
3546 => "000000000000000000000000",
3547 => "000000000000000000000000",
3548 => "000000000000000000000000",
3549 => "000000000000000000000000",
3550 => "000000000000000000000000",
3551 => "000000000000000000000000",
3552 => "000000000000000000000000",
3553 => "000000000000000000000000",
3554 => "000000000000000000000000",
3555 => "000000000000000000000000",
3556 => "000000000000000000000000",
3557 => "000000000000000000000000",
3558 => "000000000000000000000000",
3559 => "000000000000000000000000",
3560 => "000000000000000000000000",
3561 => "000000000000000000000000",
3562 => "000000000000000000000000",
3563 => "000000000000000000000000",
3564 => "000000000000000000000000",
3565 => "000000000000000000000000",
3566 => "000000000000000000000000",
3567 => "000000000000000000000000",
3568 => "000000000000000000000000",
3569 => "000000000000000000000000",
3570 => "000000000000000000000000",
3571 => "000000000000000000000000",
3572 => "000000000000000000000000",
3573 => "000000000000000000000000",
3574 => "000000000000000000000000",
3575 => "000000000000000000000000",
3576 => "000000000000000000000000",
3577 => "000000000000000000000000",
3578 => "000000000000000000000000",
3579 => "000000000000000000000000",
3580 => "000000000000000000000000",
3581 => "000000000000000000000000",
3582 => "000000000000000000000000",
3583 => "000000000000000000000000",
3584 => "000000000000000000000000",
3585 => "000000000000000000000000",
3586 => "000000000000000000000000",
3587 => "000000000000000000000000",
3588 => "000000000000000000000000",
3589 => "000000000000000000000000",
3590 => "000000000000000000000000",
3591 => "000000000000000000000000",
3592 => "000000000000000000000000",
3593 => "000000000000000000000000",
3594 => "000000000000000000000000",
3595 => "000000000000000000000000",
3596 => "000000000000000000000000",
3597 => "000000000000000000000000",
3598 => "000000000000000000000000",
3599 => "000000000000000000000000",
3600 => "000000000000000000000000",
3601 => "000000000000000000000000",
3602 => "000000000000000000000000",
3603 => "000000000000000000000000",
3604 => "000000000000000000000000",
3605 => "000000000000000000000000",
3606 => "000000000000000000000000",
3607 => "000000000000000000000000",
3608 => "000000000000000000000000",
3609 => "000000000000000000000000",
3610 => "000000000000000000000000",
3611 => "000000000000000000000000",
3612 => "000000000000000000000000",
3613 => "000000000000000000000000",
3614 => "000000000000000000000000",
3615 => "000000000000000000000000",
3616 => "000000000000000000000000",
3617 => "000000000000000000000000",
3618 => "000000000000000000000000",
3619 => "000000000000000000000000",
3620 => "000000000000000000000000",
3621 => "000000000000000000000000",
3622 => "000000000000000000000000",
3623 => "000000000000000000000000",
3624 => "000000000000000000000000",
3625 => "000000000000000000000000",
3626 => "000000000000000000000000",
3627 => "000000000000000000000000",
3628 => "000000000000000000000000",
3629 => "000000000000000000000000",
3630 => "000000000000000000000000",
3631 => "000000000000000000000000",
3632 => "000000000000000000000000",
3633 => "000000000000000000000000",
3634 => "000000000000000000000000",
3635 => "000000000000000000000000",
3636 => "000000000000000000000000",
3637 => "000000000000000000000000",
3638 => "000000000000000000000000",
3639 => "000000000000000000000000",
3640 => "000000000000000000000000",
3641 => "000000000000000000000000",
3642 => "000000000000000000000000",
3643 => "000000000000000000000000",
3644 => "000000000000000000000000",
3645 => "000000000000000000000000",
3646 => "000000000000000000000000",
3647 => "000000000000000000000000",
3648 => "000000000000000000000000",
3649 => "000000000000000000000000",
3650 => "000000000000000000000000",
3651 => "000000000000000000000000",
3652 => "000000000000000000000000",
3653 => "000000000000000000000000",
3654 => "000000000000000000000000",
3655 => "000000000000000000000000",
3656 => "000000000000000000000000",
3657 => "000000000000000000000000",
3658 => "000000000000000000000000",
3659 => "000000000000000000000000",
3660 => "000000000000000000000000",
3661 => "000000000000000000000000",
3662 => "000000000000000000000000",
3663 => "000000000000000000000000",
3664 => "000000000000000000000000",
3665 => "000110010001100100011001",
3666 => "010000110100001101000011",
3667 => "010000110100001101000011",
3668 => "010000110100001101000011",
3669 => "010000110100001101000011",
3670 => "010000110100001101000011",
3671 => "010000110100001101000011",
3672 => "001011000010110000101100",
3673 => "000000000000000000000000",
3674 => "000000000000000000000000",
3675 => "000000000000000000000000",
3676 => "000000000000000000000000",
3677 => "000000000000000000000000",
3678 => "000000000000000000000000",
3679 => "000000000000000000000000",
3680 => "000000000000000000000000",
3681 => "000000000000000000000000",
3682 => "000000000000000000000000",
3683 => "000000000000000000000000",
3684 => "000000000000000000000000",
3685 => "000000000000000000000000",
3686 => "000000000000000000000000",
3687 => "000000000000000000000000",
3688 => "000000000000000000000000",
3689 => "000000000000000000000000",
3690 => "000000000000000000000000",
3691 => "000000000000000000000000",
3692 => "000000000000000000000000",
3693 => "000000000000000000000000",
3694 => "000000000000000000000000",
3695 => "000000000000000000000000",
3696 => "000000000000000000000000",
3697 => "000000000000000000000000",
3698 => "000000000000000000000000",
3699 => "000000000000000000000000",
3700 => "000000000000000000000000",
3701 => "000000000000000000000000",
3702 => "000000000000000000000000",
3703 => "000000000000000000000000",
3704 => "000000000000000000000000",
3705 => "000000000000000000000000",
3706 => "000000000000000000000000",
3707 => "000000000000000000000000",
3708 => "000000000000000000000000",
3709 => "000000000000000000000000",
3710 => "000000000000000000000000",
3711 => "000000000000000000000000",
3712 => "000000000000000000000000",
3713 => "000000000000000000000000",
3714 => "000000000000000000000000",
3715 => "000000000000000000000000",
3716 => "000000000000000000000000",
3717 => "000000000000000000000000",
3718 => "000000000000000000000000",
3719 => "000000000000000000000000",
3720 => "000000000000000000000000",
3721 => "000000000000000000000000",
3722 => "000000000000000000000000",
3723 => "000000000000000000000000",
3724 => "000000000000000000000000",
3725 => "000000000000000000000000",
3726 => "000000000000000000000000",
3727 => "000000000000000000000000",
3728 => "000000000000000000000000",
3729 => "000000000000000000000000",
3730 => "000000000000000000000000",
3731 => "000000000000000000000000",
3732 => "000000000000000000000000",
3733 => "000000000000000000000000",
3734 => "000000000000000000000000",
3735 => "000000000000000000000000",
3736 => "000000000000000000000000",
3737 => "000000000000000000000000",
3738 => "000000000000000000000000",
3739 => "000000000000000000000000",
3740 => "000000000000000000000000",
3741 => "000000000000000000000000",
3742 => "000000000000000000000000",
3743 => "000000000000000000000000",
3744 => "000000000000000000000000",
3745 => "000000000000000000000000",
3746 => "000000000000000000000000",
3747 => "000000000000000000000000",
3748 => "000000000000000000000000",
3749 => "000000000000000000000000",
3750 => "000000000000000000000000",
3751 => "000000000000000000000000",
3752 => "000000000000000000000000",
3753 => "000000000000000000000000",
3754 => "000000000000000000000000",
3755 => "000000000000000000000000",
3756 => "000000000000000000000000",
3757 => "000000000000000000000000",
3758 => "000000000000000000000000",
3759 => "000000000000000000000000",
3760 => "000000000000000000000000",
3761 => "000000000000000000000000",
3762 => "000000000000000000000000",
3763 => "000000000000000000000000",
3764 => "000000000000000000000000",
3765 => "000000000000000000000000",
3766 => "000000000000000000000000",
3767 => "000000000000000000000000",
3768 => "000000000000000000000000",
3769 => "000000000000000000000000",
3770 => "000000000000000000000000",
3771 => "000000000000000000000000",
3772 => "000000000000000000000000",
3773 => "000000000000000000000000",
3774 => "000000000000000000000000",
3775 => "000000000000000000000000",
3776 => "000000000000000000000000",
3777 => "000000000000000000000000",
3778 => "000000000000000000000000",
3779 => "000000000000000000000000",
3780 => "000000000000000000000000",
3781 => "000000000000000000000000",
3782 => "000000000000000000000000",
3783 => "000000000000000000000000",
3784 => "000000000000000000000000",
3785 => "000000000000000000000000",
3786 => "000000000000000000000000",
3787 => "000000000000000000000000",
3788 => "000000000000000000000000",
3789 => "000000000000000000000000",
3790 => "000000000000000000000000",
3791 => "000000000000000000000000",
3792 => "000000000000000000000000",
3793 => "000000000000000000000000",
3794 => "000000000000000000000000",
3795 => "000000000000000000000000",
3796 => "000000000000000000000000",
3797 => "000000000000000000000000",
3798 => "000000000000000000000000",
3799 => "000000000000000000000000",
3800 => "000000000000000000000000",
3801 => "000000000000000000000000",
3802 => "000000000000000000000000",
3803 => "000000000000000000000000",
3804 => "000000000000000000000000",
3805 => "000000000000000000000000",
3806 => "000000000000000000000000",
3807 => "000000000000000000000000",
3808 => "000000000000000000000000",
3809 => "000000000000000000000000",
3810 => "000000000000000000000000",
3811 => "000000000000000000000000",
3812 => "000000000000000000000000",
3813 => "000010110000101100001011",
3814 => "000011110000111100001111",
3815 => "001000100010001000100010",
3816 => "010000110100001101000011",
3817 => "010000110100001101000011",
3818 => "010000110100001101000011",
3819 => "010000110100001101000011",
3820 => "010000110100001101000011",
3821 => "010000110100001101000011",
3822 => "001100010011000100110001",
3823 => "000011110000111100001111",
3824 => "000011110000111100001111",
3825 => "000000000000000000000000",
3826 => "000000000000000000000000",
3827 => "000000000000000000000000",
3828 => "000000000000000000000000",
3829 => "000000000000000000000000",
3830 => "000000000000000000000000",
3831 => "000000000000000000000000",
3832 => "000000000000000000000000",
3833 => "000000000000000000000000",
3834 => "000000000000000000000000",
3835 => "000000000000000000000000",
3836 => "000000000000000000000000",
3837 => "000000000000000000000000",
3838 => "000000000000000000000000",
3839 => "000000000000000000000000",
3840 => "000000000000000000000000",
3841 => "000000000000000000000000",
3842 => "000000000000000000000000",
3843 => "000000000000000000000000",
3844 => "000000000000000000000000",
3845 => "000000000000000000000000",
3846 => "000000000000000000000000",
3847 => "000000000000000000000000",
3848 => "000000000000000000000000",
3849 => "000000000000000000000000",
3850 => "000000000000000000000000",
3851 => "000000000000000000000000",
3852 => "000000000000000000000000",
3853 => "000000000000000000000000",
3854 => "000000000000000000000000",
3855 => "000000000000000000000000",
3856 => "000000000000000000000000",
3857 => "000000000000000000000000",
3858 => "000000000000000000000000",
3859 => "000000000000000000000000",
3860 => "000000000000000000000000",
3861 => "000000000000000000000000",
3862 => "000000000000000000000000",
3863 => "000000000000000000000000",
3864 => "000000000000000000000000",
3865 => "000000000000000000000000",
3866 => "000000000000000000000000",
3867 => "000000000000000000000000",
3868 => "000000000000000000000000",
3869 => "000000000000000000000000",
3870 => "000000000000000000000000",
3871 => "000000000000000000000000",
3872 => "000000000000000000000000",
3873 => "000000000000000000000000",
3874 => "000000000000000000000000",
3875 => "000000000000000000000000",
3876 => "000000000000000000000000",
3877 => "000000000000000000000000",
3878 => "000000000000000000000000",
3879 => "000000000000000000000000",
3880 => "000000000000000000000000",
3881 => "000000000000000000000000",
3882 => "000000000000000000000000",
3883 => "000000000000000000000000",
3884 => "000000000000000000000000",
3885 => "000000000000000000000000",
3886 => "000000000000000000000000",
3887 => "000000000000000000000000",
3888 => "000000000000000000000000",
3889 => "000000000000000000000000",
3890 => "000000000000000000000000",
3891 => "000000000000000000000000",
3892 => "000000000000000000000000",
3893 => "000000000000000000000000",
3894 => "000000000000000000000000",
3895 => "000000000000000000000000",
3896 => "000000000000000000000000",
3897 => "000000000000000000000000",
3898 => "000000000000000000000000",
3899 => "000000000000000000000000",
3900 => "000000000000000000000000",
3901 => "000000000000000000000000",
3902 => "000000000000000000000000",
3903 => "000000000000000000000000",
3904 => "000000000000000000000000",
3905 => "000000000000000000000000",
3906 => "000000000000000000000000",
3907 => "000000000000000000000000",
3908 => "000000000000000000000000",
3909 => "000000000000000000000000",
3910 => "000000000000000000000000",
3911 => "000000000000000000000000",
3912 => "000000000000000000000000",
3913 => "000000000000000000000000",
3914 => "000000000000000000000000",
3915 => "000000000000000000000000",
3916 => "000000000000000000000000",
3917 => "000000000000000000000000",
3918 => "000000000000000000000000",
3919 => "000000000000000000000000",
3920 => "000000000000000000000000",
3921 => "000000000000000000000000",
3922 => "000000000000000000000000",
3923 => "000000000000000000000000",
3924 => "000000000000000000000000",
3925 => "000000000000000000000000",
3926 => "000000000000000000000000",
3927 => "000000000000000000000000",
3928 => "000000000000000000000000",
3929 => "000000000000000000000000",
3930 => "000000000000000000000000",
3931 => "000000000000000000000000",
3932 => "000000000000000000000000",
3933 => "000000000000000000000000",
3934 => "000000000000000000000000",
3935 => "000000000000000000000000",
3936 => "000000000000000000000000",
3937 => "000000000000000000000000",
3938 => "000000000000000000000000",
3939 => "000000000000000000000000",
3940 => "000000000000000000000000",
3941 => "000000000000000000000000",
3942 => "000000000000000000000000",
3943 => "000000000000000000000000",
3944 => "000000000000000000000000",
3945 => "000000000000000000000000",
3946 => "000000000000000000000000",
3947 => "000000000000000000000000",
3948 => "000000000000000000000000",
3949 => "000000000000000000000000",
3950 => "000000000000000000000000",
3951 => "000000000000000000000000",
3952 => "000000000000000000000000",
3953 => "000000000000000000000000",
3954 => "000000000000000000000000",
3955 => "000000000000000000000000",
3956 => "000000000000000000000000",
3957 => "000000000000000000000000",
3958 => "000000000000000000000000",
3959 => "000000000000000000000000",
3960 => "000000000000000000000000",
3961 => "000000000000000000000000",
3962 => "000000000000000000000000",
3963 => "001100010011000100110001",
3964 => "010000110100001101000011",
3965 => "010000110100001101000011",
3966 => "010000110100001101000011",
3967 => "010000110100001101000011",
3968 => "010000110100001101000011",
3969 => "010000110100001101000011",
3970 => "010000110100001101000011",
3971 => "010000110100001101000011",
3972 => "010000110100001101000011",
3973 => "010000110100001101000011",
3974 => "010000110100001101000011",
3975 => "000000000000000000000000",
3976 => "000000000000000000000000",
3977 => "000000000000000000000000",
3978 => "000000000000000000000000",
3979 => "000000000000000000000000",
3980 => "000000000000000000000000",
3981 => "000000000000000000000000",
3982 => "000000000000000000000000",
3983 => "000000000000000000000000",
3984 => "000000000000000000000000",
3985 => "000000000000000000000000",
3986 => "000000000000000000000000",
3987 => "000000000000000000000000",
3988 => "000000000000000000000000",
3989 => "000000000000000000000000",
3990 => "000000000000000000000000",
3991 => "000000000000000000000000",
3992 => "000000000000000000000000",
3993 => "000000000000000000000000",
3994 => "000000000000000000000000",
3995 => "000000000000000000000000",
3996 => "000000000000000000000000",
3997 => "000000000000000000000000",
3998 => "000000000000000000000000",
3999 => "000000000000000000000000",
4000 => "000000000000000000000000",
4001 => "000000000000000000000000",
4002 => "000000000000000000000000",
4003 => "000000000000000000000000",
4004 => "000000000000000000000000",
4005 => "000000000000000000000000",
4006 => "000000000000000000000000",
4007 => "000000000000000000000000",
4008 => "000000000000000000000000",
4009 => "000000000000000000000000",
4010 => "000000000000000000000000",
4011 => "000000000000000000000000",
4012 => "000000000000000000000000",
4013 => "000000000000000000000000",
4014 => "000000000000000000000000",
4015 => "000000000000000000000000",
4016 => "000000000000000000000000",
4017 => "000000000000000000000000",
4018 => "000000000000000000000000",
4019 => "000000000000000000000000",
4020 => "000000000000000000000000",
4021 => "000000000000000000000000",
4022 => "000000000000000000000000",
4023 => "000000000000000000000000",
4024 => "000000000000000000000000",
4025 => "000000000000000000000000",
4026 => "000000000000000000000000",
4027 => "000000000000000000000000",
4028 => "000000000000000000000000",
4029 => "000000000000000000000000",
4030 => "000000000000000000000000",
4031 => "000000000000000000000000",
4032 => "000000000000000000000000",
4033 => "000000000000000000000000",
4034 => "000000000000000000000000",
4035 => "000000000000000000000000",
4036 => "000000000000000000000000",
4037 => "000000000000000000000000",
4038 => "000000000000000000000000",
4039 => "000000000000000000000000",
4040 => "000000000000000000000000",
4041 => "000000000000000000000000",
4042 => "000000000000000000000000",
4043 => "000000000000000000000000",
4044 => "000000000000000000000000",
4045 => "000000000000000000000000",
4046 => "000000000000000000000000",
4047 => "000000000000000000000000",
4048 => "000000000000000000000000",
4049 => "000000000000000000000000",
4050 => "000000000000000000000000",
4051 => "000000000000000000000000",
4052 => "000000000000000000000000",
4053 => "000000000000000000000000",
4054 => "000000000000000000000000",
4055 => "000000000000000000000000",
4056 => "000000000000000000000000",
4057 => "000000000000000000000000",
4058 => "000000000000000000000000",
4059 => "000000000000000000000000",
4060 => "000000000000000000000000",
4061 => "000000000000000000000000",
4062 => "000000000000000000000000",
4063 => "000000000000000000000000",
4064 => "000000000000000000000000",
4065 => "000000000000000000000000",
4066 => "000000000000000000000000",
4067 => "000000000000000000000000",
4068 => "000000000000000000000000",
4069 => "000000000000000000000000",
4070 => "000000000000000000000000",
4071 => "000000000000000000000000",
4072 => "000000000000000000000000",
4073 => "000000000000000000000000",
4074 => "000000000000000000000000",
4075 => "000000000000000000000000",
4076 => "000000000000000000000000",
4077 => "000000000000000000000000",
4078 => "000000000000000000000000",
4079 => "000000000000000000000000",
4080 => "000000000000000000000000",
4081 => "000000000000000000000000",
4082 => "000000000000000000000000",
4083 => "000000000000000000000000",
4084 => "000000000000000000000000",
4085 => "000000000000000000000000",
4086 => "000000000000000000000000",
4087 => "000000000000000000000000",
4088 => "000000000000000000000000",
4089 => "000000000000000000000000",
4090 => "000000000000000000000000",
4091 => "000000000000000000000000",
4092 => "000000000000000000000000",
4093 => "000000000000000000000000",
4094 => "000000000000000000000000",
4095 => "000000000000000000000000",
4096 => "000000000000000000000000",
4097 => "000000000000000000000000",
4098 => "000000000000000000000000",
4099 => "000000000000000000000000",
4100 => "000000000000000000000000",
4101 => "000000000000000000000000",
4102 => "000000000000000000000000",
4103 => "000000000000000000000000",
4104 => "000000000000000000000000",
4105 => "000000000000000000000000",
4106 => "000000000000000000000000",
4107 => "000000000000000000000000",
4108 => "000000000000000000000000",
4109 => "000000000000000000000000",
4110 => "000000000000000000000000",
4111 => "000000000000000000000000",
4112 => "000000000000000000000000",
4113 => "001100010011000100110001",
4114 => "010000110100001101000011",
4115 => "010000110100001101000011",
4116 => "010000110100001101000011",
4117 => "010000110100001101000011",
4118 => "010000110100001101000011",
4119 => "010000110100001101000011",
4120 => "010000110100001101000011",
4121 => "010000110100001101000011",
4122 => "010000110100001101000011",
4123 => "010000110100001101000011",
4124 => "010000110100001101000011",
4125 => "000000000000000000000000",
4126 => "000000000000000000000000",
4127 => "000000000000000000000000",
4128 => "000000000000000000000000",
4129 => "000000000000000000000000",
4130 => "000000000000000000000000",
4131 => "000000000000000000000000",
4132 => "000000000000000000000000",
4133 => "000000000000000000000000",
4134 => "000000000000000000000000",
4135 => "000000000000000000000000",
4136 => "000000000000000000000000",
4137 => "000000000000000000000000",
4138 => "000000000000000000000000",
4139 => "000000000000000000000000",
4140 => "000000000000000000000000",
4141 => "000000000000000000000000",
4142 => "000000000000000000000000",
4143 => "000000000000000000000000",
4144 => "000000000000000000000000",
4145 => "000000000000000000000000",
4146 => "000000000000000000000000",
4147 => "000000000000000000000000",
4148 => "000000000000000000000000",
4149 => "000000000000000000000000",
4150 => "000000000000000000000000",
4151 => "000000000000000000000000",
4152 => "000000000000000000000000",
4153 => "000000000000000000000000",
4154 => "000000000000000000000000",
4155 => "000000000000000000000000",
4156 => "000000000000000000000000",
4157 => "000000000000000000000000",
4158 => "000000000000000000000000",
4159 => "000000000000000000000000",
4160 => "000000000000000000000000",
4161 => "000000000000000000000000",
4162 => "000000000000000000000000",
4163 => "000000000000000000000000",
4164 => "000000000000000000000000",
4165 => "000000000000000000000000",
4166 => "000000000000000000000000",
4167 => "000000000000000000000000",
4168 => "000000000000000000000000",
4169 => "000000000000000000000000",
4170 => "000000000000000000000000",
4171 => "000000000000000000000000",
4172 => "000000000000000000000000",
4173 => "000000000000000000000000",
4174 => "000000000000000000000000",
4175 => "000000000000000000000000",
4176 => "000000000000000000000000",
4177 => "000000000000000000000000",
4178 => "000000000000000000000000",
4179 => "000000000000000000000000",
4180 => "000000000000000000000000",
4181 => "000000000000000000000000",
4182 => "000000000000000000000000",
4183 => "000000000000000000000000",
4184 => "000000000000000000000000",
4185 => "000000000000000000000000",
4186 => "000000000000000000000000",
4187 => "000000000000000000000000",
4188 => "000000000000000000000000",
4189 => "000000000000000000000000",
4190 => "000000000000000000000000",
4191 => "000000000000000000000000",
4192 => "000000000000000000000000",
4193 => "000000000000000000000000",
4194 => "000000000000000000000000",
4195 => "000000000000000000000000",
4196 => "000000000000000000000000",
4197 => "000000000000000000000000",
4198 => "000000000000000000000000",
4199 => "000000000000000000000000",
4200 => "000000000000000000000000",
4201 => "000000000000000000000000",
4202 => "000000000000000000000000",
4203 => "000000000000000000000000",
4204 => "000000000000000000000000",
4205 => "000000000000000000000000",
4206 => "000000000000000000000000",
4207 => "000000000000000000000000",
4208 => "000000000000000000000000",
4209 => "000000000000000000000000",
4210 => "000000000000000000000000",
4211 => "000000000000000000000000",
4212 => "000000000000000000000000",
4213 => "000000000000000000000000",
4214 => "000000000000000000000000",
4215 => "000000000000000000000000",
4216 => "000000000000000000000000",
4217 => "000000000000000000000000",
4218 => "000000000000000000000000",
4219 => "000000000000000000000000",
4220 => "000000000000000000000000",
4221 => "000000000000000000000000",
4222 => "000000000000000000000000",
4223 => "000000000000000000000000",
4224 => "000000000000000000000000",
4225 => "000000000000000000000000",
4226 => "000000000000000000000000",
4227 => "000000000000000000000000",
4228 => "000000000000000000000000",
4229 => "000000000000000000000000",
4230 => "000000000000000000000000",
4231 => "000000000000000000000000",
4232 => "000000000000000000000000",
4233 => "000000000000000000000000",
4234 => "000000000000000000000000",
4235 => "000000000000000000000000",
4236 => "000000000000000000000000",
4237 => "000000000000000000000000",
4238 => "000000000000000000000000",
4239 => "000000000000000000000000",
4240 => "000000000000000000000000",
4241 => "000000000000000000000000",
4242 => "000000000000000000000000",
4243 => "000000000000000000000000",
4244 => "000000000000000000000000",
4245 => "000000000000000000000000",
4246 => "000000000000000000000000",
4247 => "000000000000000000000000",
4248 => "000000000000000000000000",
4249 => "000000000000000000000000",
4250 => "000000000000000000000000",
4251 => "000000000000000000000000",
4252 => "000000000000000000000000",
4253 => "000000000000000000000000",
4254 => "000000000000000000000000",
4255 => "000000000000000000000000",
4256 => "000000000000000000000000",
4257 => "000000000000000000000000",
4258 => "000000000000000000000000",
4259 => "000000000000000000000000",
4260 => "000000000000000000000000",
4261 => "000000000000000000000000",
4262 => "000000000000000000000000",
4263 => "001100010011000100110001",
4264 => "010000110100001101000011",
4265 => "010000110100001101000011",
4266 => "010000110100001101000011",
4267 => "010000010100000101000001",
4268 => "000001000000010000000100",
4269 => "000001000000010000000100",
4270 => "001011110010111100101111",
4271 => "010000110100001101000011",
4272 => "010000110100001101000011",
4273 => "010000110100001101000011",
4274 => "010000110100001101000011",
4275 => "000000000000000000000000",
4276 => "000000000000000000000000",
4277 => "000000000000000000000000",
4278 => "000000000000000000000000",
4279 => "000000000000000000000000",
4280 => "000000000000000000000000",
4281 => "000000000000000000000000",
4282 => "000000000000000000000000",
4283 => "000000000000000000000000",
4284 => "000000000000000000000000",
4285 => "000000000000000000000000",
4286 => "000000000000000000000000",
4287 => "000000000000000000000000",
4288 => "000000000000000000000000",
4289 => "000000000000000000000000",
4290 => "000000000000000000000000",
4291 => "000000000000000000000000",
4292 => "000000000000000000000000",
4293 => "000000000000000000000000",
4294 => "000000000000000000000000",
4295 => "000000000000000000000000",
4296 => "000000000000000000000000",
4297 => "000000000000000000000000",
4298 => "000000000000000000000000",
4299 => "000000000000000000000000",
4300 => "000000000000000000000000",
4301 => "000000000000000000000000",
4302 => "000000000000000000000000",
4303 => "000000000000000000000000",
4304 => "000000000000000000000000",
4305 => "000000000000000000000000",
4306 => "000000000000000000000000",
4307 => "000000000000000000000000",
4308 => "000000000000000000000000",
4309 => "000000000000000000000000",
4310 => "000000000000000000000000",
4311 => "000000000000000000000000",
4312 => "000000000000000000000000",
4313 => "000000000000000000000000",
4314 => "000000000000000000000000",
4315 => "000000000000000000000000",
4316 => "000000000000000000000000",
4317 => "000000000000000000000000",
4318 => "000000000000000000000000",
4319 => "000000000000000000000000",
4320 => "000000000000000000000000",
4321 => "000000000000000000000000",
4322 => "000000000000000000000000",
4323 => "000000000000000000000000",
4324 => "000000000000000000000000",
4325 => "000000000000000000000000",
4326 => "000000000000000000000000",
4327 => "000000000000000000000000",
4328 => "000000000000000000000000",
4329 => "000000000000000000000000",
4330 => "000000000000000000000000",
4331 => "000000000000000000000000",
4332 => "000000000000000000000000",
4333 => "000000000000000000000000",
4334 => "000000000000000000000000",
4335 => "000000000000000000000000",
4336 => "000000000000000000000000",
4337 => "000000000000000000000000",
4338 => "000000000000000000000000",
4339 => "000000000000000000000000",
4340 => "000000000000000000000000",
4341 => "000000000000000000000000",
4342 => "000000000000000000000000",
4343 => "000000000000000000000000",
4344 => "000000000000000000000000",
4345 => "000000000000000000000000",
4346 => "000000000000000000000000",
4347 => "000000000000000000000000",
4348 => "000000000000000000000000",
4349 => "000000000000000000000000",
4350 => "000000000000000000000000",
4351 => "000000000000000000000000",
4352 => "000000000000000000000000",
4353 => "000000000000000000000000",
4354 => "000000000000000000000000",
4355 => "000000000000000000000000",
4356 => "000000000000000000000000",
4357 => "000000000000000000000000",
4358 => "000000000000000000000000",
4359 => "000000000000000000000000",
4360 => "000000000000000000000000",
4361 => "000000000000000000000000",
4362 => "000000000000000000000000",
4363 => "000000000000000000000000",
4364 => "000000000000000000000000",
4365 => "000000000000000000000000",
4366 => "000000000000000000000000",
4367 => "000000000000000000000000",
4368 => "000000000000000000000000",
4369 => "000000000000000000000000",
4370 => "000000000000000000000000",
4371 => "000000000000000000000000",
4372 => "000000000000000000000000",
4373 => "000000000000000000000000",
4374 => "000000000000000000000000",
4375 => "000000000000000000000000",
4376 => "000000000000000000000000",
4377 => "000000000000000000000000",
4378 => "000000000000000000000000",
4379 => "000000000000000000000000",
4380 => "000000000000000000000000",
4381 => "000000000000000000000000",
4382 => "000000000000000000000000",
4383 => "000000000000000000000000",
4384 => "000000000000000000000000",
4385 => "000000000000000000000000",
4386 => "000000000000000000000000",
4387 => "000000000000000000000000",
4388 => "000000000000000000000000",
4389 => "000000000000000000000000",
4390 => "000000000000000000000000",
4391 => "000000000000000000000000",
4392 => "000000000000000000000000",
4393 => "000000000000000000000000",
4394 => "000000000000000000000000",
4395 => "000000000000000000000000",
4396 => "000000000000000000000000",
4397 => "000000000000000000000000",
4398 => "000000000000000000000000",
4399 => "000000000000000000000000",
4400 => "000000000000000000000000",
4401 => "000000000000000000000000",
4402 => "000000000000000000000000",
4403 => "000000000000000000000000",
4404 => "000000000000000000000000",
4405 => "000000000000000000000000",
4406 => "000000000000000000000000",
4407 => "000000000000000000000000",
4408 => "000000000000000000000000",
4409 => "000000000000000000000000",
4410 => "000000000000000000000000",
4411 => "000000000000000000000000",
4412 => "000000000000000000000000",
4413 => "001100010011000100110001",
4414 => "010000110100001101000011",
4415 => "010000110100001101000011",
4416 => "010000110100001101000011",
4417 => "010000010100000101000001",
4418 => "000000000000000000000000",
4419 => "000000000000000000000000",
4420 => "001011100010111000101110",
4421 => "010000110100001101000011",
4422 => "010000110100001101000011",
4423 => "010000110100001101000011",
4424 => "010000110100001101000011",
4425 => "000000000000000000000000",
4426 => "000000000000000000000000",
4427 => "000000000000000000000000",
4428 => "000000000000000000000000",
4429 => "000000000000000000000000",
4430 => "000000000000000000000000",
4431 => "000000000000000000000000",
4432 => "000000000000000000000000",
4433 => "000000000000000000000000",
4434 => "000000000000000000000000",
4435 => "000000000000000000000000",
4436 => "000000000000000000000000",
4437 => "000000000000000000000000",
4438 => "000000000000000000000000",
4439 => "000000000000000000000000",
4440 => "000000000000000000000000",
4441 => "000000000000000000000000",
4442 => "000000000000000000000000",
4443 => "000000000000000000000000",
4444 => "000000000000000000000000",
4445 => "000000000000000000000000",
4446 => "000000000000000000000000",
4447 => "000000000000000000000000",
4448 => "000000000000000000000000",
4449 => "000000000000000000000000",
4450 => "000000000000000000000000",
4451 => "000000000000000000000000",
4452 => "000000000000000000000000",
4453 => "000000000000000000000000",
4454 => "000000000000000000000000",
4455 => "000000000000000000000000",
4456 => "000000000000000000000000",
4457 => "000000000000000000000000",
4458 => "000000000000000000000000",
4459 => "000000000000000000000000",
4460 => "000000000000000000000000",
4461 => "000000000000000000000000",
4462 => "000000000000000000000000",
4463 => "000000000000000000000000",
4464 => "000000000000000000000000",
4465 => "000000000000000000000000",
4466 => "000000000000000000000000",
4467 => "000000000000000000000000",
4468 => "000000000000000000000000",
4469 => "000000000000000000000000",
4470 => "000000000000000000000000",
4471 => "000000000000000000000000",
4472 => "000000000000000000000000",
4473 => "000000000000000000000000",
4474 => "000000000000000000000000",
4475 => "000000000000000000000000",
4476 => "000000000000000000000000",
4477 => "000000000000000000000000",
4478 => "000000000000000000000000",
4479 => "000000000000000000000000",
4480 => "000000000000000000000000",
4481 => "000000000000000000000000",
4482 => "000000000000000000000000",
4483 => "000000000000000000000000",
4484 => "000000000000000000000000",
4485 => "000000000000000000000000",
4486 => "000000000000000000000000",
4487 => "000000000000000000000000",
4488 => "000000000000000000000000",
4489 => "000000000000000000000000",
4490 => "000000000000000000000000",
4491 => "000000000000000000000000",
4492 => "000000000000000000000000",
4493 => "000000000000000000000000",
4494 => "000000000000000000000000",
4495 => "000000000000000000000000",
4496 => "000000000000000000000000",
4497 => "000000000000000000000000",
4498 => "000000000000000000000000",
4499 => "000000000000000000000000",
4500 => "000000000000000000000000",
4501 => "000000000000000000000000",
4502 => "000000000000000000000000",
4503 => "000000000000000000000000",
4504 => "000000000000000000000000",
4505 => "000000000000000000000000",
4506 => "000000000000000000000000",
4507 => "000000000000000000000000",
4508 => "000000000000000000000000",
4509 => "000000000000000000000000",
4510 => "000000000000000000000000",
4511 => "000000000000000000000000",
4512 => "000000000000000000000000",
4513 => "000000000000000000000000",
4514 => "000000000000000000000000",
4515 => "000000000000000000000000",
4516 => "000000000000000000000000",
4517 => "000000000000000000000000",
4518 => "000000000000000000000000",
4519 => "000000000000000000000000",
4520 => "000000000000000000000000",
4521 => "000000000000000000000000",
4522 => "000000000000000000000000",
4523 => "000000000000000000000000",
4524 => "000000000000000000000000",
4525 => "000000000000000000000000",
4526 => "000000000000000000000000",
4527 => "000000000000000000000000",
4528 => "000000000000000000000000",
4529 => "000000000000000000000000",
4530 => "000000000000000000000000",
4531 => "000000000000000000000000",
4532 => "000000000000000000000000",
4533 => "000000000000000000000000",
4534 => "000000000000000000000000",
4535 => "000000000000000000000000",
4536 => "000000000000000000000000",
4537 => "000000000000000000000000",
4538 => "000000000000000000000000",
4539 => "000000000000000000000000",
4540 => "000000000000000000000000",
4541 => "000000000000000000000000",
4542 => "000000000000000000000000",
4543 => "000000000000000000000000",
4544 => "000000000000000000000000",
4545 => "000000000000000000000000",
4546 => "000000000000000000000000",
4547 => "000000000000000000000000",
4548 => "000000000000000000000000",
4549 => "000000000000000000000000",
4550 => "000000000000000000000000",
4551 => "000000000000000000000000",
4552 => "000000000000000000000000",
4553 => "000000000000000000000000",
4554 => "000000000000000000000000",
4555 => "000000000000000000000000",
4556 => "000000000000000000000000",
4557 => "000000000000000000000000",
4558 => "000000000000000000000000",
4559 => "000000000000000000000000",
4560 => "000000000000000000000000",
4561 => "000000000000000000000000",
4562 => "000000000000000000000000",
4563 => "001100010011000100110001",
4564 => "010000110100001101000011",
4565 => "001101100011011000110110",
4566 => "000111110001111100011111",
4567 => "001000010010001000100010",
4568 => "010101000110100101111011",
4569 => "010101000110100101111011",
4570 => "001100000011011000111100",
4571 => "000111110001111100011111",
4572 => "001011000010110000101100",
4573 => "010000110100001101000011",
4574 => "010000110100001101000011",
4575 => "000000000000000000000000",
4576 => "000000000000000000000000",
4577 => "000000000000000000000000",
4578 => "000000000000000000000000",
4579 => "000000000000000000000000",
4580 => "000000000000000000000000",
4581 => "000000000000000000000000",
4582 => "000000000000000000000000",
4583 => "000000000000000000000000",
4584 => "000000000000000000000000",
4585 => "000000000000000000000000",
4586 => "000000000000000000000000",
4587 => "000000000000000000000000",
4588 => "000000000000000000000000",
4589 => "000000000000000000000000",
4590 => "000000000000000000000000",
4591 => "000000000000000000000000",
4592 => "000000000000000000000000",
4593 => "000000000000000000000000",
4594 => "000000000000000000000000",
4595 => "000000000000000000000000",
4596 => "000000000000000000000000",
4597 => "000000000000000000000000",
4598 => "000000000000000000000000",
4599 => "000000000000000000000000",
4600 => "000000000000000000000000",
4601 => "000000000000000000000000",
4602 => "000000000000000000000000",
4603 => "000000000000000000000000",
4604 => "000000000000000000000000",
4605 => "000000000000000000000000",
4606 => "000000000000000000000000",
4607 => "000000000000000000000000",
4608 => "000000000000000000000000",
4609 => "000000000000000000000000",
4610 => "000000000000000000000000",
4611 => "000000000000000000000000",
4612 => "000000000000000000000000",
4613 => "000000000000000000000000",
4614 => "000000000000000000000000",
4615 => "000000000000000000000000",
4616 => "000000000000000000000000",
4617 => "000000000000000000000000",
4618 => "000000000000000000000000",
4619 => "000000000000000000000000",
4620 => "000000000000000000000000",
4621 => "000000000000000000000000",
4622 => "000000000000000000000000",
4623 => "000000000000000000000000",
4624 => "000000000000000000000000",
4625 => "000000000000000000000000",
4626 => "000000000000000000000000",
4627 => "000000000000000000000000",
4628 => "000000000000000000000000",
4629 => "000000000000000000000000",
4630 => "000000000000000000000000",
4631 => "000000000000000000000000",
4632 => "000000000000000000000000",
4633 => "000000000000000000000000",
4634 => "000000000000000000000000",
4635 => "000000000000000000000000",
4636 => "000000000000000000000000",
4637 => "000000000000000000000000",
4638 => "000000000000000000000000",
4639 => "000000000000000000000000",
4640 => "000000000000000000000000",
4641 => "000000000000000000000000",
4642 => "000000000000000000000000",
4643 => "000000000000000000000000",
4644 => "000000000000000000000000",
4645 => "000000000000000000000000",
4646 => "000000000000000000000000",
4647 => "000000000000000000000000",
4648 => "000000000000000000000000",
4649 => "000000000000000000000000",
4650 => "000000000000000000000000",
4651 => "000000000000000000000000",
4652 => "000000000000000000000000",
4653 => "000000000000000000000000",
4654 => "000000000000000000000000",
4655 => "000000000000000000000000",
4656 => "000000000000000000000000",
4657 => "000000000000000000000000",
4658 => "000000000000000000000000",
4659 => "000000000000000000000000",
4660 => "000000000000000000000000",
4661 => "000000000000000000000000",
4662 => "000000000000000000000000",
4663 => "000000000000000000000000",
4664 => "000000000000000000000000",
4665 => "000000000000000000000000",
4666 => "000000000000000000000000",
4667 => "000000000000000000000000",
4668 => "000000000000000000000000",
4669 => "000000000000000000000000",
4670 => "000000000000000000000000",
4671 => "000000000000000000000000",
4672 => "000000000000000000000000",
4673 => "000000000000000000000000",
4674 => "000000000000000000000000",
4675 => "000000000000000000000000",
4676 => "000000000000000000000000",
4677 => "000000000000000000000000",
4678 => "000000000000000000000000",
4679 => "000000000000000000000000",
4680 => "000000000000000000000000",
4681 => "000000000000000000000000",
4682 => "000000000000000000000000",
4683 => "000000000000000000000000",
4684 => "000000000000000000000000",
4685 => "000000000000000000000000",
4686 => "000000000000000000000000",
4687 => "000000000000000000000000",
4688 => "000000000000000000000000",
4689 => "000000000000000000000000",
4690 => "000000000000000000000000",
4691 => "000000000000000000000000",
4692 => "000000000000000000000000",
4693 => "000000000000000000000000",
4694 => "000000000000000000000000",
4695 => "000000000000000000000000",
4696 => "000000000000000000000000",
4697 => "000000000000000000000000",
4698 => "000000000000000000000000",
4699 => "000000000000000000000000",
4700 => "000000000000000000000000",
4701 => "000000000000000000000000",
4702 => "000000000000000000000000",
4703 => "000000000000000000000000",
4704 => "000000000000000000000000",
4705 => "000000000000000000000000",
4706 => "000000000000000000000000",
4707 => "000000000000000000000000",
4708 => "000000000000000000000000",
4709 => "000000000000000000000000",
4710 => "000000000000000000000000",
4711 => "000000000000000000000000",
4712 => "000000000000000000000000",
4713 => "001100010011000100110001",
4714 => "010000110100001101000011",
4715 => "001010100010101000101010",
4716 => "000000000000000000000000",
4717 => "000001010000011000000111",
4718 => "100111111100010111101000",
4719 => "100111111100010111101000",
4720 => "001100100011111001001001",
4721 => "000000000000000000000000",
4722 => "000101110001011100010111",
4723 => "010000110100001101000011",
4724 => "010000110100001101000011",
4725 => "000000000000000000000000",
4726 => "000000000000000000000000",
4727 => "000000000000000000000000",
4728 => "000000000000000000000000",
4729 => "000000000000000000000000",
4730 => "000000000000000000000000",
4731 => "000000000000000000000000",
4732 => "000000000000000000000000",
4733 => "000000000000000000000000",
4734 => "000000000000000000000000",
4735 => "000000000000000000000000",
4736 => "000000000000000000000000",
4737 => "000000000000000000000000",
4738 => "000000000000000000000000",
4739 => "000000000000000000000000",
4740 => "000000000000000000000000",
4741 => "000000000000000000000000",
4742 => "000000000000000000000000",
4743 => "000000000000000000000000",
4744 => "000000000000000000000000",
4745 => "000000000000000000000000",
4746 => "000000000000000000000000",
4747 => "000000000000000000000000",
4748 => "000000000000000000000000",
4749 => "000000000000000000000000",
4750 => "000000000000000000000000",
4751 => "000000000000000000000000",
4752 => "000000000000000000000000",
4753 => "000000000000000000000000",
4754 => "000000000000000000000000",
4755 => "000000000000000000000000",
4756 => "000000000000000000000000",
4757 => "000000000000000000000000",
4758 => "000000000000000000000000",
4759 => "000000000000000000000000",
4760 => "000000000000000000000000",
4761 => "000000000000000000000000",
4762 => "000000000000000000000000",
4763 => "000000000000000000000000",
4764 => "000000000000000000000000",
4765 => "000000000000000000000000",
4766 => "000000000000000000000000",
4767 => "000000000000000000000000",
4768 => "000000000000000000000000",
4769 => "000000000000000000000000",
4770 => "000000000000000000000000",
4771 => "000000000000000000000000",
4772 => "000000000000000000000000",
4773 => "000000000000000000000000",
4774 => "000000000000000000000000",
4775 => "000000000000000000000000",
4776 => "000000000000000000000000",
4777 => "000000000000000000000000",
4778 => "000000000000000000000000",
4779 => "000000000000000000000000",
4780 => "000000000000000000000000",
4781 => "000000000000000000000000",
4782 => "000000000000000000000000",
4783 => "000000000000000000000000",
4784 => "000000000000000000000000",
4785 => "000000000000000000000000",
4786 => "000000000000000000000000",
4787 => "000000000000000000000000",
4788 => "000000000000000000000000",
4789 => "000000000000000000000000",
4790 => "000000000000000000000000",
4791 => "000000000000000000000000",
4792 => "000000000000000000000000",
4793 => "000000000000000000000000",
4794 => "000000000000000000000000",
4795 => "000000000000000000000000",
4796 => "000000000000000000000000",
4797 => "000000000000000000000000",
4798 => "000000000000000000000000",
4799 => "000000000000000000000000",
4800 => "000000000000000000000000",
4801 => "000000000000000000000000",
4802 => "000000000000000000000000",
4803 => "000000000000000000000000",
4804 => "000000000000000000000000",
4805 => "000000000000000000000000",
4806 => "000000000000000000000000",
4807 => "000000000000000000000000",
4808 => "000000000000000000000000",
4809 => "000000000000000000000000",
4810 => "000000000000000000000000",
4811 => "000000000000000000000000",
4812 => "000000000000000000000000",
4813 => "000000000000000000000000",
4814 => "000000000000000000000000",
4815 => "000000000000000000000000",
4816 => "000000000000000000000000",
4817 => "000000000000000000000000",
4818 => "000000000000000000000000",
4819 => "000000000000000000000000",
4820 => "000000000000000000000000",
4821 => "000000000000000000000000",
4822 => "000000000000000000000000",
4823 => "000000000000000000000000",
4824 => "000000000000000000000000",
4825 => "000000000000000000000000",
4826 => "000000000000000000000000",
4827 => "000000000000000000000000",
4828 => "000000000000000000000000",
4829 => "000000000000000000000000",
4830 => "000000000000000000000000",
4831 => "000000000000000000000000",
4832 => "000000000000000000000000",
4833 => "000000000000000000000000",
4834 => "000000000000000000000000",
4835 => "000000000000000000000000",
4836 => "000000000000000000000000",
4837 => "000000000000000000000000",
4838 => "000000000000000000000000",
4839 => "000000000000000000000000",
4840 => "000000000000000000000000",
4841 => "000000000000000000000000",
4842 => "000000000000000000000000",
4843 => "000000000000000000000000",
4844 => "000000000000000000000000",
4845 => "000000000000000000000000",
4846 => "000000000000000000000000",
4847 => "000000000000000000000000",
4848 => "000000000000000000000000",
4849 => "000000000000000000000000",
4850 => "000000000000000000000000",
4851 => "000000000000000000000000",
4852 => "000000000000000000000000",
4853 => "000000000000000000000000",
4854 => "000000000000000000000000",
4855 => "000000000000000000000000",
4856 => "000000000000000000000000",
4857 => "000000000000000000000000",
4858 => "000000000000000000000000",
4859 => "000000000000000000000000",
4860 => "000000000000000000000000",
4861 => "000000000000000000000000",
4862 => "000000000000000000000000",
4863 => "001100010011000100110001",
4864 => "010000110100001101000011",
4865 => "001010100010101000101010",
4866 => "000000000000000000000000",
4867 => "000001010000011000000111",
4868 => "100111111100010111101000",
4869 => "100111111100010111101000",
4870 => "001100100011111001001001",
4871 => "000000000000000000000000",
4872 => "000101110001011100010111",
4873 => "010000110100001101000011",
4874 => "010000110100001101000011",
4875 => "000000000000000000000000",
4876 => "000000000000000000000000",
4877 => "000000000000000000000000",
4878 => "000000000000000000000000",
4879 => "000000000000000000000000",
4880 => "000000000000000000000000",
4881 => "000000000000000000000000",
4882 => "000000000000000000000000",
4883 => "000000000000000000000000",
4884 => "000000000000000000000000",
4885 => "000000000000000000000000",
4886 => "000000000000000000000000",
4887 => "000000000000000000000000",
4888 => "000000000000000000000000",
4889 => "000000000000000000000000",
4890 => "000000000000000000000000",
4891 => "000000000000000000000000",
4892 => "000000000000000000000000",
4893 => "000000000000000000000000",
4894 => "000000000000000000000000",
4895 => "000000000000000000000000",
4896 => "000000000000000000000000",
4897 => "000000000000000000000000",
4898 => "000000000000000000000000",
4899 => "000000000000000000000000",
4900 => "000000000000000000000000",
4901 => "000000000000000000000000",
4902 => "000000000000000000000000",
4903 => "000000000000000000000000",
4904 => "000000000000000000000000",
4905 => "000000000000000000000000",
4906 => "000000000000000000000000",
4907 => "000000000000000000000000",
4908 => "000000000000000000000000",
4909 => "000000000000000000000000",
4910 => "000000000000000000000000",
4911 => "000000000000000000000000",
4912 => "000000000000000000000000",
4913 => "000000000000000000000000",
4914 => "000000000000000000000000",
4915 => "000000000000000000000000",
4916 => "000000000000000000000000",
4917 => "000000000000000000000000",
4918 => "000000000000000000000000",
4919 => "000000000000000000000000",
4920 => "000000000000000000000000",
4921 => "000000000000000000000000",
4922 => "000000000000000000000000",
4923 => "000000000000000000000000",
4924 => "000000000000000000000000",
4925 => "000000000000000000000000",
4926 => "000000000000000000000000",
4927 => "000000000000000000000000",
4928 => "000000000000000000000000",
4929 => "000000000000000000000000",
4930 => "000000000000000000000000",
4931 => "000000000000000000000000",
4932 => "000000000000000000000000",
4933 => "000000000000000000000000",
4934 => "000000000000000000000000",
4935 => "000000000000000000000000",
4936 => "000000000000000000000000",
4937 => "000000000000000000000000",
4938 => "000000000000000000000000",
4939 => "000000000000000000000000",
4940 => "000000000000000000000000",
4941 => "000000000000000000000000",
4942 => "000000000000000000000000",
4943 => "000000000000000000000000",
4944 => "000000000000000000000000",
4945 => "000000000000000000000000",
4946 => "000000000000000000000000",
4947 => "000000000000000000000000",
4948 => "000000000000000000000000",
4949 => "000000000000000000000000",
4950 => "000000000000000000000000",
4951 => "000000000000000000000000",
4952 => "000000000000000000000000",
4953 => "000000000000000000000000",
4954 => "000000000000000000000000",
4955 => "000000000000000000000000",
4956 => "000000000000000000000000",
4957 => "000000000000000000000000",
4958 => "000000000000000000000000",
4959 => "000000000000000000000000",
4960 => "000000000000000000000000",
4961 => "000000000000000000000000",
4962 => "000000000000000000000000",
4963 => "000000000000000000000000",
4964 => "000000000000000000000000",
4965 => "000000000000000000000000",
4966 => "000000000000000000000000",
4967 => "000000000000000000000000",
4968 => "000000000000000000000000",
4969 => "000000000000000000000000",
4970 => "000000000000000000000000",
4971 => "000000000000000000000000",
4972 => "000000000000000000000000",
4973 => "000000000000000000000000",
4974 => "000000000000000000000000",
4975 => "000000000000000000000000",
4976 => "000000000000000000000000",
4977 => "000000000000000000000000",
4978 => "000000000000000000000000",
4979 => "000000000000000000000000",
4980 => "000000000000000000000000",
4981 => "000000000000000000000000",
4982 => "000000000000000000000000",
4983 => "000000000000000000000000",
4984 => "000000000000000000000000",
4985 => "000000000000000000000000",
4986 => "000000000000000000000000",
4987 => "000000000000000000000000",
4988 => "000000000000000000000000",
4989 => "000000000000000000000000",
4990 => "000000000000000000000000",
4991 => "000000000000000000000000",
4992 => "000000000000000000000000",
4993 => "000000000000000000000000",
4994 => "000000000000000000000000",
4995 => "000000000000000000000000",
4996 => "000000000000000000000000",
4997 => "000000000000000000000000",
4998 => "000000000000000000000000",
4999 => "000000000000000000000000",
5000 => "000000000000000000000000",
5001 => "000000000000000000000000",
5002 => "000000000000000000000000",
5003 => "000000000000000000000000",
5004 => "000000000000000000000000",
5005 => "000000000000000000000000",
5006 => "000000000000000000000000",
5007 => "000000000000000000000000",
5008 => "000000000000000000000000",
5009 => "000000000000000000000000",
5010 => "000000000000000000000000",
5011 => "000000000000000000000000",
5012 => "000000000000000000000000",
5013 => "001100010011000100110001",
5014 => "010000110100001101000011",
5015 => "001010100010101000101010",
5016 => "000000000000000000000000",
5017 => "000001010000011000000111",
5018 => "100111111100010111101000",
5019 => "100111111100010111101000",
5020 => "001100100011111001001001",
5021 => "000000000000000000000000",
5022 => "000101110001011100010111",
5023 => "010000110100001101000011",
5024 => "010000110100001101000011",
5025 => "000000000000000000000000",
5026 => "000000000000000000000000",
5027 => "000000000000000000000000",
5028 => "000000000000000000000000",
5029 => "000000000000000000000000",
5030 => "000000000000000000000000",
5031 => "000000000000000000000000",
5032 => "000000000000000000000000",
5033 => "000000000000000000000000",
5034 => "000000000000000000000000",
5035 => "000000000000000000000000",
5036 => "000000000000000000000000",
5037 => "000000000000000000000000",
5038 => "000000000000000000000000",
5039 => "000000000000000000000000",
5040 => "000000000000000000000000",
5041 => "000000000000000000000000",
5042 => "000000000000000000000000",
5043 => "000000000000000000000000",
5044 => "000000000000000000000000",
5045 => "000000000000000000000000",
5046 => "000000000000000000000000",
5047 => "000000000000000000000000",
5048 => "000000000000000000000000",
5049 => "000000000000000000000000",
5050 => "000000000000000000000000",
5051 => "000000000000000000000000",
5052 => "000000000000000000000000",
5053 => "000000000000000000000000",
5054 => "000000000000000000000000",
5055 => "000000000000000000000000",
5056 => "000000000000000000000000",
5057 => "000000000000000000000000",
5058 => "000000000000000000000000",
5059 => "000000000000000000000000",
5060 => "000000000000000000000000",
5061 => "000000000000000000000000",
5062 => "000000000000000000000000",
5063 => "000000000000000000000000",
5064 => "000000000000000000000000",
5065 => "000000000000000000000000",
5066 => "000000000000000000000000",
5067 => "000000000000000000000000",
5068 => "000000000000000000000000",
5069 => "000000000000000000000000",
5070 => "000000000000000000000000",
5071 => "000000000000000000000000",
5072 => "000000000000000000000000",
5073 => "000000000000000000000000",
5074 => "000000000000000000000000",
5075 => "000000000000000000000000",
5076 => "000000000000000000000000",
5077 => "000000000000000000000000",
5078 => "000000000000000000000000",
5079 => "000000000000000000000000",
5080 => "000000000000000000000000",
5081 => "000000000000000000000000",
5082 => "000000000000000000000000",
5083 => "000000000000000000000000",
5084 => "000000000000000000000000",
5085 => "000000000000000000000000",
5086 => "000000000000000000000000",
5087 => "000000000000000000000000",
5088 => "000000000000000000000000",
5089 => "000000000000000000000000",
5090 => "000000000000000000000000",
5091 => "000000000000000000000000",
5092 => "000000000000000000000000",
5093 => "000000000000000000000000",
5094 => "000000000000000000000000",
5095 => "000000000000000000000000",
5096 => "000000000000000000000000",
5097 => "000000000000000000000000",
5098 => "000000000000000000000000",
5099 => "000000000000000000000000",
5100 => "000000000000000000000000",
5101 => "000000000000000000000000",
5102 => "000000000000000000000000",
5103 => "000000000000000000000000",
5104 => "000000000000000000000000",
5105 => "000000000000000000000000",
5106 => "000000000000000000000000",
5107 => "000000000000000000000000",
5108 => "000000000000000000000000",
5109 => "000000000000000000000000",
5110 => "000000000000000000000000",
5111 => "000000000000000000000000",
5112 => "000000000000000000000000",
5113 => "000000000000000000000000",
5114 => "000000000000000000000000",
5115 => "000000000000000000000000",
5116 => "000000000000000000000000",
5117 => "000000000000000000000000",
5118 => "000000000000000000000000",
5119 => "000000000000000000000000",
5120 => "000000000000000000000000",
5121 => "000000000000000000000000",
5122 => "000000000000000000000000",
5123 => "000000000000000000000000",
5124 => "000000000000000000000000",
5125 => "000000000000000000000000",
5126 => "000000000000000000000000",
5127 => "000000000000000000000000",
5128 => "000000000000000000000000",
5129 => "000000000000000000000000",
5130 => "000000000000000000000000",
5131 => "000000000000000000000000",
5132 => "000000000000000000000000",
5133 => "000000000000000000000000",
5134 => "000000000000000000000000",
5135 => "000000000000000000000000",
5136 => "000000000000000000000000",
5137 => "000000000000000000000000",
5138 => "000000000000000000000000",
5139 => "000000000000000000000000",
5140 => "000000000000000000000000",
5141 => "000000000000000000000000",
5142 => "000000000000000000000000",
5143 => "000000000000000000000000",
5144 => "000000000000000000000000",
5145 => "000000000000000000000000",
5146 => "000000000000000000000000",
5147 => "000000000000000000000000",
5148 => "000000000000000000000000",
5149 => "000000000000000000000000",
5150 => "000000000000000000000000",
5151 => "000000000000000000000000",
5152 => "000000000000000000000000",
5153 => "000000000000000000000000",
5154 => "000000000000000000000000",
5155 => "000000000000000000000000",
5156 => "000000000000000000000000",
5157 => "000000000000000000000000",
5158 => "000000000000000000000000",
5159 => "000000000000000000000000",
5160 => "000000000000000000000000",
5161 => "000000000000000000000000",
5162 => "000000000000000000000000",
5163 => "001100010011000100110001",
5164 => "010000110100001101000011",
5165 => "001010100010101000101010",
5166 => "000000000000000000000000",
5167 => "000001010000011000000111",
5168 => "100111111100010111101000",
5169 => "100111111100010111101000",
5170 => "001100100011111001001001",
5171 => "000000000000000000000000",
5172 => "000101110001011100010111",
5173 => "010000110100001101000011",
5174 => "010000110100001101000011",
5175 => "000000000000000000000000",
5176 => "000000000000000000000000",
5177 => "000000000000000000000000",
5178 => "000000000000000000000000",
5179 => "000000000000000000000000",
5180 => "000000000000000000000000",
5181 => "000000000000000000000000",
5182 => "000000000000000000000000",
5183 => "000000000000000000000000",
5184 => "000000000000000000000000",
5185 => "000000000000000000000000",
5186 => "000000000000000000000000",
5187 => "000000000000000000000000",
5188 => "000000000000000000000000",
5189 => "000000000000000000000000",
5190 => "000000000000000000000000",
5191 => "000000000000000000000000",
5192 => "000000000000000000000000",
5193 => "000000000000000000000000",
5194 => "000000000000000000000000",
5195 => "000000000000000000000000",
5196 => "000000000000000000000000",
5197 => "000000000000000000000000",
5198 => "000000000000000000000000",
5199 => "000000000000000000000000",
5200 => "000000000000000000000000",
5201 => "000000000000000000000000",
5202 => "000000000000000000000000",
5203 => "000000000000000000000000",
5204 => "000000000000000000000000",
5205 => "000000000000000000000000",
5206 => "000000000000000000000000",
5207 => "000000000000000000000000",
5208 => "000000000000000000000000",
5209 => "000000000000000000000000",
5210 => "000000000000000000000000",
5211 => "000000000000000000000000",
5212 => "000000000000000000000000",
5213 => "000000000000000000000000",
5214 => "000000000000000000000000",
5215 => "000000000000000000000000",
5216 => "000000000000000000000000",
5217 => "000000000000000000000000",
5218 => "000000000000000000000000",
5219 => "000000000000000000000000",
5220 => "000000000000000000000000",
5221 => "000000000000000000000000",
5222 => "000000000000000000000000",
5223 => "000000000000000000000000",
5224 => "000000000000000000000000",
5225 => "000000000000000000000000",
5226 => "000000000000000000000000",
5227 => "000000000000000000000000",
5228 => "000000000000000000000000",
5229 => "000000000000000000000000",
5230 => "000000000000000000000000",
5231 => "000000000000000000000000",
5232 => "000000000000000000000000",
5233 => "000000000000000000000000",
5234 => "000000000000000000000000",
5235 => "000000000000000000000000",
5236 => "000000000000000000000000",
5237 => "000000000000000000000000",
5238 => "000000000000000000000000",
5239 => "000000000000000000000000",
5240 => "000000000000000000000000",
5241 => "000000000000000000000000",
5242 => "000000000000000000000000",
5243 => "000000000000000000000000",
5244 => "000000000000000000000000",
5245 => "000000000000000000000000",
5246 => "000000000000000000000000",
5247 => "000000000000000000000000",
5248 => "000000000000000000000000",
5249 => "000000000000000000000000",
5250 => "000000000000000000000000",
5251 => "000000000000000000000000",
5252 => "000000000000000000000000",
5253 => "000000000000000000000000",
5254 => "000000000000000000000000",
5255 => "000000000000000000000000",
5256 => "000000000000000000000000",
5257 => "000000000000000000000000",
5258 => "000000000000000000000000",
5259 => "000000000000000000000000",
5260 => "000000000000000000000000",
5261 => "000000000000000000000000",
5262 => "000000000000000000000000",
5263 => "000000000000000000000000",
5264 => "000000000000000000000000",
5265 => "000000000000000000000000",
5266 => "000000000000000000000000",
5267 => "000000000000000000000000",
5268 => "000000000000000000000000",
5269 => "000000000000000000000000",
5270 => "000000000000000000000000",
5271 => "000000000000000000000000",
5272 => "000000000000000000000000",
5273 => "000000000000000000000000",
5274 => "000000000000000000000000",
5275 => "000000000000000000000000",
5276 => "000000000000000000000000",
5277 => "000000000000000000000000",
5278 => "000000000000000000000000",
5279 => "000000000000000000000000",
5280 => "000000000000000000000000",
5281 => "000000000000000000000000",
5282 => "000000000000000000000000",
5283 => "000000000000000000000000",
5284 => "000000000000000000000000",
5285 => "000000000000000000000000",
5286 => "000000000000000000000000",
5287 => "000000000000000000000000",
5288 => "000000000000000000000000",
5289 => "000000000000000000000000",
5290 => "000000000000000000000000",
5291 => "000000000000000000000000",
5292 => "000000000000000000000000",
5293 => "000000000000000000000000",
5294 => "000000000000000000000000",
5295 => "000000000000000000000000",
5296 => "000000000000000000000000",
5297 => "000000000000000000000000",
5298 => "000000000000000000000000",
5299 => "000000000000000000000000",
5300 => "000000000000000000000000",
5301 => "000000000000000000000000",
5302 => "000000000000000000000000",
5303 => "000000000000000000000000",
5304 => "000000000000000000000000",
5305 => "000000000000000000000000",
5306 => "000000000000000000000000",
5307 => "000000000000000000000000",
5308 => "000000000000000000000000",
5309 => "000000000000000000000000",
5310 => "000001000000010000000100",
5311 => "001111010011110100111101",
5312 => "001111010011110100111101",
5313 => "000101010001010100010101",
5314 => "000001100000011000000110",
5315 => "001110100100011101010011",
5316 => "100100101011010111010101",
5317 => "100100101011010111010101",
5318 => "100111111100010111101000",
5319 => "100111111100010111101000",
5320 => "100101101011101011011011",
5321 => "100100101011010111010101",
5322 => "011000100111100010001101",
5323 => "000001100000011000000110",
5324 => "000001100000011000000110",
5325 => "001111010011110100111101",
5326 => "001111010011110100111101",
5327 => "000101010001010100010101",
5328 => "000000000000000000000000",
5329 => "000000000000000000000000",
5330 => "000000000000000000000000",
5331 => "000000000000000000000000",
5332 => "000000000000000000000000",
5333 => "000000000000000000000000",
5334 => "000000000000000000000000",
5335 => "000000000000000000000000",
5336 => "000000000000000000000000",
5337 => "000000000000000000000000",
5338 => "000000000000000000000000",
5339 => "000000000000000000000000",
5340 => "000000000000000000000000",
5341 => "000000000000000000000000",
5342 => "000000000000000000000000",
5343 => "000000000000000000000000",
5344 => "000000000000000000000000",
5345 => "000000000000000000000000",
5346 => "000000000000000000000000",
5347 => "000000000000000000000000",
5348 => "000000000000000000000000",
5349 => "000000000000000000000000",
5350 => "000000000000000000000000",
5351 => "000000000000000000000000",
5352 => "000000000000000000000000",
5353 => "000000000000000000000000",
5354 => "000000000000000000000000",
5355 => "000000000000000000000000",
5356 => "000000000000000000000000",
5357 => "000000000000000000000000",
5358 => "000000000000000000000000",
5359 => "000000000000000000000000",
5360 => "000000000000000000000000",
5361 => "000000000000000000000000",
5362 => "000000000000000000000000",
5363 => "000000000000000000000000",
5364 => "000000000000000000000000",
5365 => "000000000000000000000000",
5366 => "000000000000000000000000",
5367 => "000000000000000000000000",
5368 => "000000000000000000000000",
5369 => "000000000000000000000000",
5370 => "000000000000000000000000",
5371 => "000000000000000000000000",
5372 => "000000000000000000000000",
5373 => "000000000000000000000000",
5374 => "000000000000000000000000",
5375 => "000000000000000000000000",
5376 => "000000000000000000000000",
5377 => "000000000000000000000000",
5378 => "000000000000000000000000",
5379 => "000000000000000000000000",
5380 => "000000000000000000000000",
5381 => "000000000000000000000000",
5382 => "000000000000000000000000",
5383 => "000000000000000000000000",
5384 => "000000000000000000000000",
5385 => "000000000000000000000000",
5386 => "000000000000000000000000",
5387 => "000000000000000000000000",
5388 => "000000000000000000000000",
5389 => "000000000000000000000000",
5390 => "000000000000000000000000",
5391 => "000000000000000000000000",
5392 => "000000000000000000000000",
5393 => "000000000000000000000000",
5394 => "000000000000000000000000",
5395 => "000000000000000000000000",
5396 => "000000000000000000000000",
5397 => "000000000000000000000000",
5398 => "000000000000000000000000",
5399 => "000000000000000000000000",
5400 => "000000000000000000000000",
5401 => "000000000000000000000000",
5402 => "000000000000000000000000",
5403 => "000000000000000000000000",
5404 => "000000000000000000000000",
5405 => "000000000000000000000000",
5406 => "000000000000000000000000",
5407 => "000000000000000000000000",
5408 => "000000000000000000000000",
5409 => "000000000000000000000000",
5410 => "000000000000000000000000",
5411 => "000000000000000000000000",
5412 => "000000000000000000000000",
5413 => "000000000000000000000000",
5414 => "000000000000000000000000",
5415 => "000000000000000000000000",
5416 => "000000000000000000000000",
5417 => "000000000000000000000000",
5418 => "000000000000000000000000",
5419 => "000000000000000000000000",
5420 => "000000000000000000000000",
5421 => "000000000000000000000000",
5422 => "000000000000000000000000",
5423 => "000000000000000000000000",
5424 => "000000000000000000000000",
5425 => "000000000000000000000000",
5426 => "000000000000000000000000",
5427 => "000000000000000000000000",
5428 => "000000000000000000000000",
5429 => "000000000000000000000000",
5430 => "000000000000000000000000",
5431 => "000000000000000000000000",
5432 => "000000000000000000000000",
5433 => "000000000000000000000000",
5434 => "000000000000000000000000",
5435 => "000000000000000000000000",
5436 => "000000000000000000000000",
5437 => "000000000000000000000000",
5438 => "000000000000000000000000",
5439 => "000000000000000000000000",
5440 => "000000000000000000000000",
5441 => "000000000000000000000000",
5442 => "000000000000000000000000",
5443 => "000000000000000000000000",
5444 => "000000000000000000000000",
5445 => "000000000000000000000000",
5446 => "000000000000000000000000",
5447 => "000000000000000000000000",
5448 => "000000000000000000000000",
5449 => "000000000000000000000000",
5450 => "000000000000000000000000",
5451 => "000000000000000000000000",
5452 => "000000000000000000000000",
5453 => "000000000000000000000000",
5454 => "000000000000000000000000",
5455 => "000000000000000000000000",
5456 => "000000000000000000000000",
5457 => "000000000000000000000000",
5458 => "000000000000000000000000",
5459 => "000000000000000000000000",
5460 => "000001000000010000000100",
5461 => "010000110100001101000011",
5462 => "010000110100001101000011",
5463 => "000100100001001000010010",
5464 => "000000000000000000000000",
5465 => "001111000100101001010111",
5466 => "100111111100010111101000",
5467 => "100111111100010111101000",
5468 => "100111111100010111101000",
5469 => "100111111100010111101000",
5470 => "100111111100010111101000",
5471 => "100111111100010111101000",
5472 => "011010001000000110011000",
5473 => "000000000000000000000000",
5474 => "000000000000000000000000",
5475 => "010000110100001101000011",
5476 => "010000110100001101000011",
5477 => "000101110001011100010111",
5478 => "000000000000000000000000",
5479 => "000000000000000000000000",
5480 => "000000000000000000000000",
5481 => "000000000000000000000000",
5482 => "000000000000000000000000",
5483 => "000000000000000000000000",
5484 => "000000000000000000000000",
5485 => "000000000000000000000000",
5486 => "000000000000000000000000",
5487 => "000000000000000000000000",
5488 => "000000000000000000000000",
5489 => "000000000000000000000000",
5490 => "000000000000000000000000",
5491 => "000000000000000000000000",
5492 => "000000000000000000000000",
5493 => "000000000000000000000000",
5494 => "000000000000000000000000",
5495 => "000000000000000000000000",
5496 => "000000000000000000000000",
5497 => "000000000000000000000000",
5498 => "000000000000000000000000",
5499 => "000000000000000000000000",
5500 => "000000000000000000000000",
5501 => "000000000000000000000000",
5502 => "000000000000000000000000",
5503 => "000000000000000000000000",
5504 => "000000000000000000000000",
5505 => "000000000000000000000000",
5506 => "000000000000000000000000",
5507 => "000000000000000000000000",
5508 => "000000000000000000000000",
5509 => "000000000000000000000000",
5510 => "000000000000000000000000",
5511 => "000000000000000000000000",
5512 => "000000000000000000000000",
5513 => "000000000000000000000000",
5514 => "000000000000000000000000",
5515 => "000000000000000000000000",
5516 => "000000000000000000000000",
5517 => "000000000000000000000000",
5518 => "000000000000000000000000",
5519 => "000000000000000000000000",
5520 => "000000000000000000000000",
5521 => "000000000000000000000000",
5522 => "000000000000000000000000",
5523 => "000000000000000000000000",
5524 => "000000000000000000000000",
5525 => "000000000000000000000000",
5526 => "000000000000000000000000",
5527 => "000000000000000000000000",
5528 => "000000000000000000000000",
5529 => "000000000000000000000000",
5530 => "000000000000000000000000",
5531 => "000000000000000000000000",
5532 => "000000000000000000000000",
5533 => "000000000000000000000000",
5534 => "000000000000000000000000",
5535 => "000000000000000000000000",
5536 => "000000000000000000000000",
5537 => "000000000000000000000000",
5538 => "000000000000000000000000",
5539 => "000000000000000000000000",
5540 => "000000000000000000000000",
5541 => "000000000000000000000000",
5542 => "000000000000000000000000",
5543 => "000000000000000000000000",
5544 => "000000000000000000000000",
5545 => "000000000000000000000000",
5546 => "000000000000000000000000",
5547 => "000000000000000000000000",
5548 => "000000000000000000000000",
5549 => "000000000000000000000000",
5550 => "000000000000000000000000",
5551 => "000000000000000000000000",
5552 => "000000000000000000000000",
5553 => "000000000000000000000000",
5554 => "000000000000000000000000",
5555 => "000000000000000000000000",
5556 => "000000000000000000000000",
5557 => "000000000000000000000000",
5558 => "000000000000000000000000",
5559 => "000000000000000000000000",
5560 => "000000000000000000000000",
5561 => "000000000000000000000000",
5562 => "000000000000000000000000",
5563 => "000000000000000000000000",
5564 => "000000000000000000000000",
5565 => "000000000000000000000000",
5566 => "000000000000000000000000",
5567 => "000000000000000000000000",
5568 => "000000000000000000000000",
5569 => "000000000000000000000000",
5570 => "000000000000000000000000",
5571 => "000000000000000000000000",
5572 => "000000000000000000000000",
5573 => "000000000000000000000000",
5574 => "000000000000000000000000",
5575 => "000000000000000000000000",
5576 => "000000000000000000000000",
5577 => "000000000000000000000000",
5578 => "000000000000000000000000",
5579 => "000000000000000000000000",
5580 => "000000000000000000000000",
5581 => "000000000000000000000000",
5582 => "000000000000000000000000",
5583 => "000000000000000000000000",
5584 => "000000000000000000000000",
5585 => "000000000000000000000000",
5586 => "000000000000000000000000",
5587 => "000000000000000000000000",
5588 => "000000000000000000000000",
5589 => "000000000000000000000000",
5590 => "000000000000000000000000",
5591 => "000000000000000000000000",
5592 => "000000000000000000000000",
5593 => "000000000000000000000000",
5594 => "000000000000000000000000",
5595 => "000000000000000000000000",
5596 => "000000000000000000000000",
5597 => "000000000000000000000000",
5598 => "000000000000000000000000",
5599 => "000000000000000000000000",
5600 => "000000000000000000000000",
5601 => "000000000000000000000000",
5602 => "000000000000000000000000",
5603 => "000000000000000000000000",
5604 => "000000000000000000000000",
5605 => "000000000000000000000000",
5606 => "000000000000000000000000",
5607 => "000000000000000000000000",
5608 => "000000000000000000000000",
5609 => "000000000000000000000000",
5610 => "000001000000010000000100",
5611 => "010000110100001101000011",
5612 => "010000110100001101000011",
5613 => "000100100001001000010010",
5614 => "000000000000000000000000",
5615 => "001111000100101001010111",
5616 => "100111111100010111101000",
5617 => "100111111100010111101000",
5618 => "100111111100010111101000",
5619 => "100111111100010111101000",
5620 => "100111111100010111101000",
5621 => "100111111100010111101000",
5622 => "011010001000000110011000",
5623 => "000000000000000000000000",
5624 => "000000000000000000000000",
5625 => "010000110100001101000011",
5626 => "010000110100001101000011",
5627 => "000101110001011100010111",
5628 => "000000000000000000000000",
5629 => "000000000000000000000000",
5630 => "000000000000000000000000",
5631 => "000000000000000000000000",
5632 => "000000000000000000000000",
5633 => "000000000000000000000000",
5634 => "000000000000000000000000",
5635 => "000000000000000000000000",
5636 => "000000000000000000000000",
5637 => "000000000000000000000000",
5638 => "000000000000000000000000",
5639 => "000000000000000000000000",
5640 => "000000000000000000000000",
5641 => "000000000000000000000000",
5642 => "000000000000000000000000",
5643 => "000000000000000000000000",
5644 => "000000000000000000000000",
5645 => "000000000000000000000000",
5646 => "000000000000000000000000",
5647 => "000000000000000000000000",
5648 => "000000000000000000000000",
5649 => "000000000000000000000000",
5650 => "000000000000000000000000",
5651 => "000000000000000000000000",
5652 => "000000000000000000000000",
5653 => "000000000000000000000000",
5654 => "000000000000000000000000",
5655 => "000000000000000000000000",
5656 => "000000000000000000000000",
5657 => "000000000000000000000000",
5658 => "000000000000000000000000",
5659 => "000000000000000000000000",
5660 => "000000000000000000000000",
5661 => "000000000000000000000000",
5662 => "000000000000000000000000",
5663 => "000000000000000000000000",
5664 => "000000000000000000000000",
5665 => "000000000000000000000000",
5666 => "000000000000000000000000",
5667 => "000000000000000000000000",
5668 => "000000000000000000000000",
5669 => "000000000000000000000000",
5670 => "000000000000000000000000",
5671 => "000000000000000000000000",
5672 => "000000000000000000000000",
5673 => "000000000000000000000000",
5674 => "000000000000000000000000",
5675 => "000000000000000000000000",
5676 => "000000000000000000000000",
5677 => "000000000000000000000000",
5678 => "000000000000000000000000",
5679 => "000000000000000000000000",
5680 => "000000000000000000000000",
5681 => "000000000000000000000000",
5682 => "000000000000000000000000",
5683 => "000000000000000000000000",
5684 => "000000000000000000000000",
5685 => "000000000000000000000000",
5686 => "000000000000000000000000",
5687 => "000000000000000000000000",
5688 => "000000000000000000000000",
5689 => "000000000000000000000000",
5690 => "000000000000000000000000",
5691 => "000000000000000000000000",
5692 => "000000000000000000000000",
5693 => "000000000000000000000000",
5694 => "000000000000000000000000",
5695 => "000000000000000000000000",
5696 => "000000000000000000000000",
5697 => "000000000000000000000000",
5698 => "000000000000000000000000",
5699 => "000000000000000000000000",
5700 => "000000000000000000000000",
5701 => "000000000000000000000000",
5702 => "000000000000000000000000",
5703 => "000000000000000000000000",
5704 => "000000000000000000000000",
5705 => "000000000000000000000000",
5706 => "000000000000000000000000",
5707 => "000000000000000000000000",
5708 => "000000000000000000000000",
5709 => "000000000000000000000000",
5710 => "000000000000000000000000",
5711 => "000000000000000000000000",
5712 => "000000000000000000000000",
5713 => "000000000000000000000000",
5714 => "000000000000000000000000",
5715 => "000000000000000000000000",
5716 => "000000000000000000000000",
5717 => "000000000000000000000000",
5718 => "000000000000000000000000",
5719 => "000000000000000000000000",
5720 => "000000000000000000000000",
5721 => "000000000000000000000000",
5722 => "000000000000000000000000",
5723 => "000000000000000000000000",
5724 => "000000000000000000000000",
5725 => "000000000000000000000000",
5726 => "000000000000000000000000",
5727 => "000000000000000000000000",
5728 => "000000000000000000000000",
5729 => "000000000000000000000000",
5730 => "000000000000000000000000",
5731 => "000000000000000000000000",
5732 => "000000000000000000000000",
5733 => "000000000000000000000000",
5734 => "000000000000000000000000",
5735 => "000000000000000000000000",
5736 => "000000000000000000000000",
5737 => "000000000000000000000000",
5738 => "000000000000000000000000",
5739 => "000000000000000000000000",
5740 => "000000000000000000000000",
5741 => "000000000000000000000000",
5742 => "000000000000000000000000",
5743 => "000000000000000000000000",
5744 => "000000000000000000000000",
5745 => "000000000000000000000000",
5746 => "000000000000000000000000",
5747 => "000000000000000000000000",
5748 => "000000000000000000000000",
5749 => "000000000000000000000000",
5750 => "000000000000000000000000",
5751 => "000000000000000000000000",
5752 => "000000000000000000000000",
5753 => "000000000000000000000000",
5754 => "000000000000000000000000",
5755 => "000000000000000000000000",
5756 => "000000000000000000000000",
5757 => "000000000000000000000000",
5758 => "000000000000000000000000",
5759 => "000000000000000000000000",
5760 => "000001000000010000000100",
5761 => "010000110100001101000011",
5762 => "010000110100001101000011",
5763 => "000100100001001000010010",
5764 => "000000000000000000000000",
5765 => "001111000100101001010111",
5766 => "100111111100010111101000",
5767 => "100111111100010111101000",
5768 => "100111111100010111101000",
5769 => "100111111100010111101000",
5770 => "100111111100010111101000",
5771 => "100111111100010111101000",
5772 => "011010001000000110011000",
5773 => "000000000000000000000000",
5774 => "000000000000000000000000",
5775 => "010000110100001101000011",
5776 => "010000110100001101000011",
5777 => "000101110001011100010111",
5778 => "000000000000000000000000",
5779 => "000000000000000000000000",
5780 => "000000000000000000000000",
5781 => "000000000000000000000000",
5782 => "000000000000000000000000",
5783 => "000000000000000000000000",
5784 => "000000000000000000000000",
5785 => "000000000000000000000000",
5786 => "000000000000000000000000",
5787 => "000000000000000000000000",
5788 => "000000000000000000000000",
5789 => "000000000000000000000000",
5790 => "000000000000000000000000",
5791 => "000000000000000000000000",
5792 => "000000000000000000000000",
5793 => "000000000000000000000000",
5794 => "000000000000000000000000",
5795 => "000000000000000000000000",
5796 => "000000000000000000000000",
5797 => "000000000000000000000000",
5798 => "000000000000000000000000",
5799 => "000000000000000000000000",
5800 => "000000000000000000000000",
5801 => "000000000000000000000000",
5802 => "000000000000000000000000",
5803 => "000000000000000000000000",
5804 => "000000000000000000000000",
5805 => "000000000000000000000000",
5806 => "000000000000000000000000",
5807 => "000000000000000000000000",
5808 => "000000000000000000000000",
5809 => "000000000000000000000000",
5810 => "000000000000000000000000",
5811 => "000000000000000000000000",
5812 => "000000000000000000000000",
5813 => "000000000000000000000000",
5814 => "000000000000000000000000",
5815 => "000000000000000000000000",
5816 => "000000000000000000000000",
5817 => "000000000000000000000000",
5818 => "000000000000000000000000",
5819 => "000000000000000000000000",
5820 => "000000000000000000000000",
5821 => "000000000000000000000000",
5822 => "000000000000000000000000",
5823 => "000000000000000000000000",
5824 => "000000000000000000000000",
5825 => "000000000000000000000000",
5826 => "000000000000000000000000",
5827 => "000000000000000000000000",
5828 => "000000000000000000000000",
5829 => "000000000000000000000000",
5830 => "000000000000000000000000",
5831 => "000000000000000000000000",
5832 => "000000000000000000000000",
5833 => "000000000000000000000000",
5834 => "000000000000000000000000",
5835 => "000000000000000000000000",
5836 => "000000000000000000000000",
5837 => "000000000000000000000000",
5838 => "000000000000000000000000",
5839 => "000000000000000000000000",
5840 => "000000000000000000000000",
5841 => "000000000000000000000000",
5842 => "000000000000000000000000",
5843 => "000000000000000000000000",
5844 => "000000000000000000000000",
5845 => "000000000000000000000000",
5846 => "000000000000000000000000",
5847 => "000000000000000000000000",
5848 => "000000000000000000000000",
5849 => "000000000000000000000000",
5850 => "000000000000000000000000",
5851 => "000000000000000000000000",
5852 => "000000000000000000000000",
5853 => "000000000000000000000000",
5854 => "000000000000000000000000",
5855 => "000000000000000000000000",
5856 => "000000000000000000000000",
5857 => "000000000000000000000000",
5858 => "000000000000000000000000",
5859 => "000000000000000000000000",
5860 => "000000000000000000000000",
5861 => "000000000000000000000000",
5862 => "000000000000000000000000",
5863 => "000000000000000000000000",
5864 => "000000000000000000000000",
5865 => "000000000000000000000000",
5866 => "000000000000000000000000",
5867 => "000000000000000000000000",
5868 => "000000000000000000000000",
5869 => "000000000000000000000000",
5870 => "000000000000000000000000",
5871 => "000000000000000000000000",
5872 => "000000000000000000000000",
5873 => "000000000000000000000000",
5874 => "000000000000000000000000",
5875 => "000000000000000000000000",
5876 => "000000000000000000000000",
5877 => "000000000000000000000000",
5878 => "000000000000000000000000",
5879 => "000000000000000000000000",
5880 => "000000000000000000000000",
5881 => "000000000000000000000000",
5882 => "000000000000000000000000",
5883 => "000000000000000000000000",
5884 => "000000000000000000000000",
5885 => "000000000000000000000000",
5886 => "000000000000000000000000",
5887 => "000000000000000000000000",
5888 => "000000000000000000000000",
5889 => "000000000000000000000000",
5890 => "000000000000000000000000",
5891 => "000000000000000000000000",
5892 => "000000000000000000000000",
5893 => "000000000000000000000000",
5894 => "000000000000000000000000",
5895 => "000000000000000000000000",
5896 => "000000000000000000000000",
5897 => "000000000000000000000000",
5898 => "000000000000000000000000",
5899 => "000000000000000000000000",
5900 => "000000000000000000000000",
5901 => "000000000000000000000000",
5902 => "000000000000000000000000",
5903 => "000000000000000000000000",
5904 => "000000000000000000000000",
5905 => "000000000000000000000000",
5906 => "000000000000000000000000",
5907 => "000000000000000000000000",
5908 => "000000000000000000000000",
5909 => "000000000000000000000000",
5910 => "000001000000010000000100",
5911 => "010000110100001101000011",
5912 => "010000110100001101000011",
5913 => "000100100001001000010010",
5914 => "000000000000000000000000",
5915 => "001111000100101001010111",
5916 => "100111111100010111101000",
5917 => "100111111100010111101000",
5918 => "100111111100010111101000",
5919 => "100111111100010111101000",
5920 => "100111111100010111101000",
5921 => "100111111100010111101000",
5922 => "011010001000000110011000",
5923 => "000000000000000000000000",
5924 => "000000000000000000000000",
5925 => "010000110100001101000011",
5926 => "010000110100001101000011",
5927 => "000101110001011100010111",
5928 => "000000000000000000000000",
5929 => "000000000000000000000000",
5930 => "000000000000000000000000",
5931 => "000000000000000000000000",
5932 => "000000000000000000000000",
5933 => "000000000000000000000000",
5934 => "000000000000000000000000",
5935 => "000000000000000000000000",
5936 => "000000000000000000000000",
5937 => "000000000000000000000000",
5938 => "000000000000000000000000",
5939 => "000000000000000000000000",
5940 => "000000000000000000000000",
5941 => "000000000000000000000000",
5942 => "000000000000000000000000",
5943 => "000000000000000000000000",
5944 => "000000000000000000000000",
5945 => "000000000000000000000000",
5946 => "000000000000000000000000",
5947 => "000000000000000000000000",
5948 => "000000000000000000000000",
5949 => "000000000000000000000000",
5950 => "000000000000000000000000",
5951 => "000000000000000000000000",
5952 => "000000000000000000000000",
5953 => "000000000000000000000000",
5954 => "000000000000000000000000",
5955 => "000000000000000000000000",
5956 => "000000000000000000000000",
5957 => "000000000000000000000000",
5958 => "000000000000000000000000",
5959 => "000000000000000000000000",
5960 => "000000000000000000000000",
5961 => "000000000000000000000000",
5962 => "000000000000000000000000",
5963 => "000000000000000000000000",
5964 => "000000000000000000000000",
5965 => "000000000000000000000000",
5966 => "000000000000000000000000",
5967 => "000000000000000000000000",
5968 => "000000000000000000000000",
5969 => "000000000000000000000000",
5970 => "000000000000000000000000",
5971 => "000000000000000000000000",
5972 => "000000000000000000000000",
5973 => "000000000000000000000000",
5974 => "000000000000000000000000",
5975 => "000000000000000000000000",
5976 => "000000000000000000000000",
5977 => "000000000000000000000000",
5978 => "000000000000000000000000",
5979 => "000000000000000000000000",
5980 => "000000000000000000000000",
5981 => "000000000000000000000000",
5982 => "000000000000000000000000",
5983 => "000000000000000000000000",
5984 => "000000000000000000000000",
5985 => "000000000000000000000000",
5986 => "000000000000000000000000",
5987 => "000000000000000000000000",
5988 => "000000000000000000000000",
5989 => "000000000000000000000000",
5990 => "000000000000000000000000",
5991 => "000000000000000000000000",
5992 => "000000000000000000000000",
5993 => "000000000000000000000000",
5994 => "000000000000000000000000",
5995 => "000000000000000000000000",
5996 => "000000000000000000000000",
5997 => "000000000000000000000000",
5998 => "000000000000000000000000",
5999 => "000000000000000000000000",
6000 => "000000000000000000000000",
6001 => "000000000000000000000000",
6002 => "000000000000000000000000",
6003 => "000000000000000000000000",
6004 => "000000000000000000000000",
6005 => "000000000000000000000000",
6006 => "000000000000000000000000",
6007 => "000000000000000000000000",
6008 => "000000000000000000000000",
6009 => "000000000000000000000000",
6010 => "000000000000000000000000",
6011 => "000000000000000000000000",
6012 => "000000000000000000000000",
6013 => "000000000000000000000000",
6014 => "000000000000000000000000",
6015 => "000000000000000000000000",
6016 => "000000000000000000000000",
6017 => "000000000000000000000000",
6018 => "000000000000000000000000",
6019 => "000000000000000000000000",
6020 => "000000000000000000000000",
6021 => "000000000000000000000000",
6022 => "000000000000000000000000",
6023 => "000000000000000000000000",
6024 => "000000000000000000000000",
6025 => "000000000000000000000000",
6026 => "000000000000000000000000",
6027 => "000000000000000000000000",
6028 => "000000000000000000000000",
6029 => "000000000000000000000000",
6030 => "000000000000000000000000",
6031 => "000000000000000000000000",
6032 => "000000000000000000000000",
6033 => "000000000000000000000000",
6034 => "000000000000000000000000",
6035 => "000000000000000000000000",
6036 => "000000000000000000000000",
6037 => "000000000000000000000000",
6038 => "000000000000000000000000",
6039 => "000000000000000000000000",
6040 => "000000000000000000000000",
6041 => "000000000000000000000000",
6042 => "000000000000000000000000",
6043 => "000000000000000000000000",
6044 => "000000000000000000000000",
6045 => "000000000000000000000000",
6046 => "000000000000000000000000",
6047 => "000000000000000000000000",
6048 => "000000000000000000000000",
6049 => "000000000000000000000000",
6050 => "000000000000000000000000",
6051 => "000000000000000000000000",
6052 => "000000000000000000000000",
6053 => "000000000000000000000000",
6054 => "000000000000000000000000",
6055 => "000000000000000000000000",
6056 => "000000000000000000000000",
6057 => "000000000000000000000000",
6058 => "000000000000000000000000",
6059 => "000000000000000000000000",
6060 => "000001000000010000000100",
6061 => "010000110100001101000011",
6062 => "010000110100001101000011",
6063 => "000100100001001000010010",
6064 => "000000000000000000000000",
6065 => "001111000100101001010111",
6066 => "100111111100010111101000",
6067 => "100111111100010111101000",
6068 => "100111111100010111101000",
6069 => "100111111100010111101000",
6070 => "100111111100010111101000",
6071 => "100111111100010111101000",
6072 => "011010001000000110011000",
6073 => "000000000000000000000000",
6074 => "000000000000000000000000",
6075 => "010000110100001101000011",
6076 => "010000110100001101000011",
6077 => "000101110001011100010111",
6078 => "000000000000000000000000",
6079 => "000000000000000000000000",
6080 => "000000000000000000000000",
6081 => "000000000000000000000000",
6082 => "000000000000000000000000",
6083 => "000000000000000000000000",
6084 => "000000000000000000000000",
6085 => "000000000000000000000000",
6086 => "000000000000000000000000",
6087 => "000000000000000000000000",
6088 => "000000000000000000000000",
6089 => "000000000000000000000000",
6090 => "000000000000000000000000",
6091 => "000000000000000000000000",
6092 => "000000000000000000000000",
6093 => "000000000000000000000000",
6094 => "000000000000000000000000",
6095 => "000000000000000000000000",
6096 => "000000000000000000000000",
6097 => "000000000000000000000000",
6098 => "000000000000000000000000",
6099 => "000000000000000000000000",
6100 => "000000000000000000000000",
6101 => "000000000000000000000000",
6102 => "000000000000000000000000",
6103 => "000000000000000000000000",
6104 => "000000000000000000000000",
6105 => "000000000000000000000000",
6106 => "000000000000000000000000",
6107 => "000000000000000000000000",
6108 => "000000000000000000000000",
6109 => "000000000000000000000000",
6110 => "000000000000000000000000",
6111 => "000000000000000000000000",
6112 => "000000000000000000000000",
6113 => "000000000000000000000000",
6114 => "000000000000000000000000",
6115 => "000000000000000000000000",
6116 => "000000000000000000000000",
6117 => "000000000000000000000000",
6118 => "000000000000000000000000",
6119 => "000000000000000000000000",
6120 => "000000000000000000000000",
6121 => "000000000000000000000000",
6122 => "000000000000000000000000",
6123 => "000000000000000000000000",
6124 => "000000000000000000000000",
6125 => "000000000000000000000000",
6126 => "000000000000000000000000",
6127 => "000000000000000000000000",
6128 => "000000000000000000000000",
6129 => "000000000000000000000000",
6130 => "000000000000000000000000",
6131 => "000000000000000000000000",
6132 => "000000000000000000000000",
6133 => "000000000000000000000000",
6134 => "000000000000000000000000",
6135 => "000000000000000000000000",
6136 => "000000000000000000000000",
6137 => "000000000000000000000000",
6138 => "000000000000000000000000",
6139 => "000000000000000000000000",
6140 => "000000000000000000000000",
6141 => "000000000000000000000000",
6142 => "000000000000000000000000",
6143 => "000000000000000000000000",
6144 => "000000000000000000000000",
6145 => "000000000000000000000000",
6146 => "000000000000000000000000",
6147 => "000000000000000000000000",
6148 => "000000000000000000000000",
6149 => "000000000000000000000000",
6150 => "000000000000000000000000",
6151 => "000000000000000000000000",
6152 => "000000000000000000000000",
6153 => "000000000000000000000000",
6154 => "000000000000000000000000",
6155 => "000000000000000000000000",
6156 => "000000000000000000000000",
6157 => "000000000000000000000000",
6158 => "000000000000000000000000",
6159 => "000000000000000000000000",
6160 => "000000000000000000000000",
6161 => "000000000000000000000000",
6162 => "000000000000000000000000",
6163 => "000000000000000000000000",
6164 => "000000000000000000000000",
6165 => "000000000000000000000000",
6166 => "000000000000000000000000",
6167 => "000000000000000000000000",
6168 => "000000000000000000000000",
6169 => "000000000000000000000000",
6170 => "000000000000000000000000",
6171 => "000000000000000000000000",
6172 => "000000000000000000000000",
6173 => "000000000000000000000000",
6174 => "000000000000000000000000",
6175 => "000000000000000000000000",
6176 => "000000000000000000000000",
6177 => "000000000000000000000000",
6178 => "000000000000000000000000",
6179 => "000000000000000000000000",
6180 => "000000000000000000000000",
6181 => "000000000000000000000000",
6182 => "000000000000000000000000",
6183 => "000000000000000000000000",
6184 => "000000000000000000000000",
6185 => "000000000000000000000000",
6186 => "000000000000000000000000",
6187 => "000000000000000000000000",
6188 => "000000000000000000000000",
6189 => "000000000000000000000000",
6190 => "000000000000000000000000",
6191 => "000000000000000000000000",
6192 => "000000000000000000000000",
6193 => "000000000000000000000000",
6194 => "000000000000000000000000",
6195 => "000000000000000000000000",
6196 => "000000000000000000000000",
6197 => "000000000000000000000000",
6198 => "000000000000000000000000",
6199 => "000000000000000000000000",
6200 => "000000000000000000000000",
6201 => "000000000000000000000000",
6202 => "000000000000000000000000",
6203 => "000000000000000000000000",
6204 => "000000000000000000000000",
6205 => "000000000000000000000000",
6206 => "000000000000000000000000",
6207 => "000000000000000000000000",
6208 => "000000000000000000000000",
6209 => "000000000000000000000000",
6210 => "000001000000010000000100",
6211 => "010000110100001101000011",
6212 => "010000110100001101000011",
6213 => "000100100001001000010010",
6214 => "000000000000000000000000",
6215 => "001111000100101001010111",
6216 => "100111111100010111101000",
6217 => "100111111100010111101000",
6218 => "100111111100010111101000",
6219 => "100111111100010111101000",
6220 => "100111111100010111101000",
6221 => "100111111100010111101000",
6222 => "011010001000000110011000",
6223 => "000000000000000000000000",
6224 => "000000000000000000000000",
6225 => "010000110100001101000011",
6226 => "010000110100001101000011",
6227 => "000101110001011100010111",
6228 => "000000000000000000000000",
6229 => "000000000000000000000000",
6230 => "000000000000000000000000",
6231 => "000000000000000000000000",
6232 => "000000000000000000000000",
6233 => "000000000000000000000000",
6234 => "000000000000000000000000",
6235 => "000000000000000000000000",
6236 => "000000000000000000000000",
6237 => "000000000000000000000000",
6238 => "000000000000000000000000",
6239 => "000000000000000000000000",
6240 => "000000000000000000000000",
6241 => "000000000000000000000000",
6242 => "000000000000000000000000",
6243 => "000000000000000000000000",
6244 => "000000000000000000000000",
6245 => "000000000000000000000000",
6246 => "000000000000000000000000",
6247 => "000000000000000000000000",
6248 => "000000000000000000000000",
6249 => "000000000000000000000000",
6250 => "000000000000000000000000",
6251 => "000000000000000000000000",
6252 => "000000000000000000000000",
6253 => "000000000000000000000000",
6254 => "000000000000000000000000",
6255 => "000000000000000000000000",
6256 => "000000000000000000000000",
6257 => "000000000000000000000000",
6258 => "000000000000000000000000",
6259 => "000000000000000000000000",
6260 => "000000000000000000000000",
6261 => "000000000000000000000000",
6262 => "000000000000000000000000",
6263 => "000000000000000000000000",
6264 => "000000000000000000000000",
6265 => "000000000000000000000000",
6266 => "000000000000000000000000",
6267 => "000000000000000000000000",
6268 => "000000000000000000000000",
6269 => "000000000000000000000000",
6270 => "000000000000000000000000",
6271 => "000000000000000000000000",
6272 => "000000000000000000000000",
6273 => "000000000000000000000000",
6274 => "000000000000000000000000",
6275 => "000000000000000000000000",
6276 => "000000000000000000000000",
6277 => "000000000000000000000000",
6278 => "000000000000000000000000",
6279 => "000000000000000000000000",
6280 => "000000000000000000000000",
6281 => "000000000000000000000000",
6282 => "000000000000000000000000",
6283 => "000000000000000000000000",
6284 => "000000000000000000000000",
6285 => "000000000000000000000000",
6286 => "000000000000000000000000",
6287 => "000000000000000000000000",
6288 => "000000000000000000000000",
6289 => "000000000000000000000000",
6290 => "000000000000000000000000",
6291 => "000000000000000000000000",
6292 => "000000000000000000000000",
6293 => "000000000000000000000000",
6294 => "000000000000000000000000",
6295 => "000000000000000000000000",
6296 => "000000000000000000000000",
6297 => "000000000000000000000000",
6298 => "000000000000000000000000",
6299 => "000000000000000000000000",
6300 => "000000000000000000000000",
6301 => "000000000000000000000000",
6302 => "000000000000000000000000",
6303 => "000000000000000000000000",
6304 => "000000000000000000000000",
6305 => "000000000000000000000000",
6306 => "000000000000000000000000",
6307 => "000000000000000000000000",
6308 => "000000000000000000000000",
6309 => "000000000000000000000000",
6310 => "000000000000000000000000",
6311 => "000000000000000000000000",
6312 => "000000000000000000000000",
6313 => "000000000000000000000000",
6314 => "000000000000000000000000",
6315 => "000000000000000000000000",
6316 => "000000000000000000000000",
6317 => "000000000000000000000000",
6318 => "000000000000000000000000",
6319 => "000000000000000000000000",
6320 => "000000000000000000000000",
6321 => "000000000000000000000000",
6322 => "000000000000000000000000",
6323 => "000000000000000000000000",
6324 => "000000000000000000000000",
6325 => "000000000000000000000000",
6326 => "000000000000000000000000",
6327 => "000000000000000000000000",
6328 => "000000000000000000000000",
6329 => "000000000000000000000000",
6330 => "000000000000000000000000",
6331 => "000000000000000000000000",
6332 => "000000000000000000000000",
6333 => "000000000000000000000000",
6334 => "000000000000000000000000",
6335 => "000000000000000000000000",
6336 => "000000000000000000000000",
6337 => "000000000000000000000000",
6338 => "000000000000000000000000",
6339 => "000000000000000000000000",
6340 => "000000000000000000000000",
6341 => "000000000000000000000000",
6342 => "000000000000000000000000",
6343 => "000000000000000000000000",
6344 => "000000000000000000000000",
6345 => "000000000000000000000000",
6346 => "000000000000000000000000",
6347 => "000000000000000000000000",
6348 => "000000000000000000000000",
6349 => "000000000000000000000000",
6350 => "000000000000000000000000",
6351 => "000000000000000000000000",
6352 => "000000000000000000000000",
6353 => "000000000000000000000000",
6354 => "000000000000000000000000",
6355 => "000000000000000000000000",
6356 => "000000000000000000000000",
6357 => "000000000000000000000000",
6358 => "000000000000000000000000",
6359 => "000000000000000000000000",
6360 => "000001000000010000000100",
6361 => "010000110100001101000011",
6362 => "010000110100001101000011",
6363 => "000100100001001000010010",
6364 => "000000000000000000000000",
6365 => "001111000100101001010111",
6366 => "100111111100010111101000",
6367 => "100111111100010111101000",
6368 => "100111111100010111101000",
6369 => "100111111100010111101000",
6370 => "100111111100010111101000",
6371 => "100111111100010111101000",
6372 => "011010001000000110011000",
6373 => "000000000000000000000000",
6374 => "000000000000000000000000",
6375 => "010000110100001101000011",
6376 => "010000110100001101000011",
6377 => "000101110001011100010111",
6378 => "000000000000000000000000",
6379 => "000000000000000000000000",
6380 => "000000000000000000000000",
6381 => "000000000000000000000000",
6382 => "000000000000000000000000",
6383 => "000000000000000000000000",
6384 => "000000000000000000000000",
6385 => "000000000000000000000000",
6386 => "000000000000000000000000",
6387 => "000000000000000000000000",
6388 => "000000000000000000000000",
6389 => "000000000000000000000000",
6390 => "000000000000000000000000",
6391 => "000000000000000000000000",
6392 => "000000000000000000000000",
6393 => "000000000000000000000000",
6394 => "000000000000000000000000",
6395 => "000000000000000000000000",
6396 => "000000000000000000000000",
6397 => "000000000000000000000000",
6398 => "000000000000000000000000",
6399 => "000000000000000000000000",
6400 => "000000000000000000000000",
6401 => "000000000000000000000000",
6402 => "000000000000000000000000",
6403 => "000000000000000000000000",
6404 => "000000000000000000000000",
6405 => "000000000000000000000000",
6406 => "000000000000000000000000",
6407 => "000000000000000000000000",
6408 => "000000000000000000000000",
6409 => "000000000000000000000000",
6410 => "000000000000000000000000",
6411 => "000000000000000000000000",
6412 => "000000000000000000000000",
6413 => "000000000000000000000000",
6414 => "000000000000000000000000",
6415 => "000000000000000000000000",
6416 => "000000000000000000000000",
6417 => "000000000000000000000000",
6418 => "000000000000000000000000",
6419 => "000000000000000000000000",
6420 => "000000000000000000000000",
6421 => "000000000000000000000000",
6422 => "000000000000000000000000",
6423 => "000000000000000000000000",
6424 => "000000000000000000000000",
6425 => "000000000000000000000000",
6426 => "000000000000000000000000",
6427 => "000000000000000000000000",
6428 => "000000000000000000000000",
6429 => "000000000000000000000000",
6430 => "000000000000000000000000",
6431 => "000000000000000000000000",
6432 => "000000000000000000000000",
6433 => "000000000000000000000000",
6434 => "000000000000000000000000",
6435 => "000000000000000000000000",
6436 => "000000000000000000000000",
6437 => "000000000000000000000000",
6438 => "000000000000000000000000",
6439 => "000000000000000000000000",
6440 => "000000000000000000000000",
6441 => "000000000000000000000000",
6442 => "000000000000000000000000",
6443 => "000000000000000000000000",
6444 => "000000000000000000000000",
6445 => "000000000000000000000000",
6446 => "000000000000000000000000",
6447 => "000000000000000000000000",
6448 => "000000000000000000000000",
6449 => "000000000000000000000000",
6450 => "000000000000000000000000",
6451 => "000000000000000000000000",
6452 => "000000000000000000000000",
6453 => "000000000000000000000000",
6454 => "000000000000000000000000",
6455 => "000000000000000000000000",
6456 => "000000000000000000000000",
6457 => "000000000000000000000000",
6458 => "000000000000000000000000",
6459 => "000000000000000000000000",
6460 => "000000000000000000000000",
6461 => "000000000000000000000000",
6462 => "000000000000000000000000",
6463 => "000000000000000000000000",
6464 => "000000000000000000000000",
6465 => "000000000000000000000000",
6466 => "000000000000000000000000",
6467 => "000000000000000000000000",
6468 => "000000000000000000000000",
6469 => "000000000000000000000000",
6470 => "000000000000000000000000",
6471 => "000000000000000000000000",
6472 => "000000000000000000000000",
6473 => "000000000000000000000000",
6474 => "000000000000000000000000",
6475 => "000000000000000000000000",
6476 => "000000000000000000000000",
6477 => "000000000000000000000000",
6478 => "000000000000000000000000",
6479 => "000000000000000000000000",
6480 => "000000000000000000000000",
6481 => "000000000000000000000000",
6482 => "000000000000000000000000",
6483 => "000000000000000000000000",
6484 => "000000000000000000000000",
6485 => "000000000000000000000000",
6486 => "000000000000000000000000",
6487 => "000000000000000000000000",
6488 => "000000000000000000000000",
6489 => "000000000000000000000000",
6490 => "000000000000000000000000",
6491 => "000000000000000000000000",
6492 => "000000000000000000000000",
6493 => "000000000000000000000000",
6494 => "000000000000000000000000",
6495 => "000000000000000000000000",
6496 => "000000000000000000000000",
6497 => "000000000000000000000000",
6498 => "000000000000000000000000",
6499 => "000000000000000000000000",
6500 => "000000000000000000000000",
6501 => "000000000000000000000000",
6502 => "000000000000000000000000",
6503 => "000000000000000000000000",
6504 => "000000000000000000000000",
6505 => "000000000000000000000000",
6506 => "000000000000000000000000",
6507 => "000000000000000000000000",
6508 => "000000000000000000000000",
6509 => "000000000000000000000000",
6510 => "000001000000010000000100",
6511 => "010000110100001101000011",
6512 => "010000110100001101000011",
6513 => "000100100001001000010010",
6514 => "000000000000000000000000",
6515 => "001111000100101001010111",
6516 => "100111111100010111101000",
6517 => "100111111100010111101000",
6518 => "100111111100010111101000",
6519 => "100111111100010111101000",
6520 => "100111111100010111101000",
6521 => "100111111100010111101000",
6522 => "011010001000000110011000",
6523 => "000000000000000000000000",
6524 => "000000000000000000000000",
6525 => "010000110100001101000011",
6526 => "010000110100001101000011",
6527 => "000101110001011100010111",
6528 => "000000000000000000000000",
6529 => "000000000000000000000000",
6530 => "000000000000000000000000",
6531 => "000000000000000000000000",
6532 => "000000000000000000000000",
6533 => "000000000000000000000000",
6534 => "000000000000000000000000",
6535 => "000000000000000000000000",
6536 => "000000000000000000000000",
6537 => "000000000000000000000000",
6538 => "000000000000000000000000",
6539 => "000000000000000000000000",
6540 => "000000000000000000000000",
6541 => "000000000000000000000000",
6542 => "000000000000000000000000",
6543 => "000000000000000000000000",
6544 => "000000000000000000000000",
6545 => "000000000000000000000000",
6546 => "000000000000000000000000",
6547 => "000000000000000000000000",
6548 => "000000000000000000000000",
6549 => "000000000000000000000000",
6550 => "000000000000000000000000",
6551 => "000000000000000000000000",
6552 => "000000000000000000000000",
6553 => "000000000000000000000000",
6554 => "000000000000000000000000",
6555 => "000000000000000000000000",
6556 => "000000000000000000000000",
6557 => "000000000000000000000000",
6558 => "000000000000000000000000",
6559 => "000000000000000000000000",
6560 => "000000000000000000000000",
6561 => "000000000000000000000000",
6562 => "000000000000000000000000",
6563 => "000000000000000000000000",
6564 => "000000000000000000000000",
6565 => "000000000000000000000000",
6566 => "000000000000000000000000",
6567 => "000000000000000000000000",
6568 => "000000000000000000000000",
6569 => "000000000000000000000000",
6570 => "000000000000000000000000",
6571 => "000000000000000000000000",
6572 => "000000000000000000000000",
6573 => "000000000000000000000000",
6574 => "000000000000000000000000",
6575 => "000000000000000000000000",
6576 => "000000000000000000000000",
6577 => "000000000000000000000000",
6578 => "000000000000000000000000",
6579 => "000000000000000000000000",
6580 => "000000000000000000000000",
6581 => "000000000000000000000000",
6582 => "000000000000000000000000",
6583 => "000000000000000000000000",
6584 => "000000000000000000000000",
6585 => "000000000000000000000000",
6586 => "000000000000000000000000",
6587 => "000000000000000000000000",
6588 => "000000000000000000000000",
6589 => "000000000000000000000000",
6590 => "000000000000000000000000",
6591 => "000000000000000000000000",
6592 => "000000000000000000000000",
6593 => "000000000000000000000000",
6594 => "000000000000000000000000",
6595 => "000000000000000000000000",
6596 => "000000000000000000000000",
6597 => "000000000000000000000000",
6598 => "000000000000000000000000",
6599 => "000000000000000000000000",
6600 => "000000000000000000000000",
6601 => "000000000000000000000000",
6602 => "000000000000000000000000",
6603 => "000000000000000000000000",
6604 => "000000000000000000000000",
6605 => "000000000000000000000000",
6606 => "000000000000000000000000",
6607 => "000000000000000000000000",
6608 => "000000000000000000000000",
6609 => "000000000000000000000000",
6610 => "000000000000000000000000",
6611 => "000000000000000000000000",
6612 => "000000000000000000000000",
6613 => "000000000000000000000000",
6614 => "000000000000000000000000",
6615 => "000000000000000000000000",
6616 => "000000000000000000000000",
6617 => "000000000000000000000000",
6618 => "000000000000000000000000",
6619 => "000000000000000000000000",
6620 => "000000000000000000000000",
6621 => "000000000000000000000000",
6622 => "000000000000000000000000",
6623 => "000000000000000000000000",
6624 => "000000000000000000000000",
6625 => "000000000000000000000000",
6626 => "000000000000000000000000",
6627 => "000000000000000000000000",
6628 => "000000000000000000000000",
6629 => "000000000000000000000000",
6630 => "000000000000000000000000",
6631 => "000000000000000000000000",
6632 => "000000000000000000000000",
6633 => "000000000000000000000000",
6634 => "000000000000000000000000",
6635 => "000000000000000000000000",
6636 => "000000000000000000000000",
6637 => "000000000000000000000000",
6638 => "000000000000000000000000",
6639 => "000000000000000000000000",
6640 => "000000000000000000000000",
6641 => "000000000000000000000000",
6642 => "000000000000000000000000",
6643 => "000000000000000000000000",
6644 => "000000000000000000000000",
6645 => "000000000000000000000000",
6646 => "000000000000000000000000",
6647 => "000000000000000000000000",
6648 => "000000000000000000000000",
6649 => "000000000000000000000000",
6650 => "000000000000000000000000",
6651 => "000000000000000000000000",
6652 => "000000000000000000000000",
6653 => "000000000000000000000000",
6654 => "000000000000000000000000",
6655 => "000000000000000000000000",
6656 => "000000000000000000000000",
6657 => "000000000000000000000000",
6658 => "000000000000000000000000",
6659 => "000000000000000000000000",
6660 => "000001000000010000000100",
6661 => "010000110100001101000011",
6662 => "010000110100001101000011",
6663 => "000100100001001000010010",
6664 => "000000000000000000000000",
6665 => "001111000100101001010111",
6666 => "100111111100010111101000",
6667 => "100111111100010111101000",
6668 => "100111111100010111101000",
6669 => "100111111100010111101000",
6670 => "100111111100010111101000",
6671 => "100111111100010111101000",
6672 => "011010001000000110011000",
6673 => "000000000000000000000000",
6674 => "000000000000000000000000",
6675 => "010000110100001101000011",
6676 => "010000110100001101000011",
6677 => "000101110001011100010111",
6678 => "000000000000000000000000",
6679 => "000000000000000000000000",
6680 => "000000000000000000000000",
6681 => "000000000000000000000000",
6682 => "000000000000000000000000",
6683 => "000000000000000000000000",
6684 => "000000000000000000000000",
6685 => "000000000000000000000000",
6686 => "000000000000000000000000",
6687 => "000000000000000000000000",
6688 => "000000000000000000000000",
6689 => "000000000000000000000000",
6690 => "000000000000000000000000",
6691 => "000000000000000000000000",
6692 => "000000000000000000000000",
6693 => "000000000000000000000000",
6694 => "000000000000000000000000",
6695 => "000000000000000000000000",
6696 => "000000000000000000000000",
6697 => "000000000000000000000000",
6698 => "000000000000000000000000",
6699 => "000000000000000000000000",
6700 => "000000000000000000000000",
6701 => "000000000000000000000000",
6702 => "000000000000000000000000",
6703 => "000000000000000000000000",
6704 => "000000000000000000000000",
6705 => "000000000000000000000000",
6706 => "000000000000000000000000",
6707 => "000000000000000000000000",
6708 => "000000000000000000000000",
6709 => "000000000000000000000000",
6710 => "000000000000000000000000",
6711 => "000000000000000000000000",
6712 => "000000000000000000000000",
6713 => "000000000000000000000000",
6714 => "000000000000000000000000",
6715 => "000000000000000000000000",
6716 => "000000000000000000000000",
6717 => "000000000000000000000000",
6718 => "000000000000000000000000",
6719 => "000000000000000000000000",
6720 => "000000000000000000000000",
6721 => "000000000000000000000000",
6722 => "000000000000000000000000",
6723 => "000000000000000000000000",
6724 => "000000000000000000000000",
6725 => "000000000000000000000000",
6726 => "000000000000000000000000",
6727 => "000000000000000000000000",
6728 => "000000000000000000000000",
6729 => "000000000000000000000000",
6730 => "000000000000000000000000",
6731 => "000000000000000000000000",
6732 => "000000000000000000000000",
6733 => "000000000000000000000000",
6734 => "000000000000000000000000",
6735 => "000000000000000000000000",
6736 => "000000000000000000000000",
6737 => "000000000000000000000000",
6738 => "000000000000000000000000",
6739 => "000000000000000000000000",
6740 => "000000000000000000000000",
6741 => "000000000000000000000000",
6742 => "000000000000000000000000",
6743 => "000000000000000000000000",
6744 => "000000000000000000000000",
6745 => "000000000000000000000000",
6746 => "000000000000000000000000",
6747 => "000000000000000000000000",
6748 => "000000000000000000000000",
6749 => "000000000000000000000000",
6750 => "000000000000000000000000",
6751 => "000000000000000000000000",
6752 => "000000000000000000000000",
6753 => "000000000000000000000000",
6754 => "000000000000000000000000",
6755 => "000000000000000000000000",
6756 => "000000000000000000000000",
6757 => "000000000000000000000000",
6758 => "000000000000000000000000",
6759 => "000000000000000000000000",
6760 => "000000000000000000000000",
6761 => "000000000000000000000000",
6762 => "000000000000000000000000",
6763 => "000000000000000000000000",
6764 => "000000000000000000000000",
6765 => "000000000000000000000000",
6766 => "000000000000000000000000",
6767 => "000000000000000000000000",
6768 => "000000000000000000000000",
6769 => "000000000000000000000000",
6770 => "000000000000000000000000",
6771 => "000000000000000000000000",
6772 => "000000000000000000000000",
6773 => "000000000000000000000000",
6774 => "000000000000000000000000",
6775 => "000000000000000000000000",
6776 => "000000000000000000000000",
6777 => "000000000000000000000000",
6778 => "000000000000000000000000",
6779 => "000000000000000000000000",
6780 => "000000000000000000000000",
6781 => "000000000000000000000000",
6782 => "000000000000000000000000",
6783 => "000000000000000000000000",
6784 => "000000000000000000000000",
6785 => "000000000000000000000000",
6786 => "000000000000000000000000",
6787 => "000000000000000000000000",
6788 => "000000000000000000000000",
6789 => "000000000000000000000000",
6790 => "000000000000000000000000",
6791 => "000000000000000000000000",
6792 => "000000000000000000000000",
6793 => "000000000000000000000000",
6794 => "000000000000000000000000",
6795 => "000000000000000000000000",
6796 => "000000000000000000000000",
6797 => "000000000000000000000000",
6798 => "000000000000000000000000",
6799 => "000000000000000000000000",
6800 => "000000000000000000000000",
6801 => "000000000000000000000000",
6802 => "000000000000000000000000",
6803 => "000000000000000000000000",
6804 => "000000000000000000000000",
6805 => "000000000000000000000000",
6806 => "000000000000000000000000",
6807 => "000000000000000000000000",
6808 => "000000000000000000000000",
6809 => "000000000000000000000000",
6810 => "000001000000010000000100",
6811 => "010000110100001101000011",
6812 => "010000110100001101000011",
6813 => "000100100001001000010010",
6814 => "000000000000000000000000",
6815 => "001111000100101001010111",
6816 => "100111111100010111101000",
6817 => "100111111100010111101000",
6818 => "100111111100010111101000",
6819 => "100111111100010111101000",
6820 => "100111111100010111101000",
6821 => "100111111100010111101000",
6822 => "011010001000000110011000",
6823 => "000000000000000000000000",
6824 => "000000000000000000000000",
6825 => "010000110100001101000011",
6826 => "010000110100001101000011",
6827 => "000101110001011100010111",
6828 => "000000000000000000000000",
6829 => "000000000000000000000000",
6830 => "000000000000000000000000",
6831 => "000000000000000000000000",
6832 => "000000000000000000000000",
6833 => "000000000000000000000000",
6834 => "000000000000000000000000",
6835 => "000000000000000000000000",
6836 => "000000000000000000000000",
6837 => "000000000000000000000000",
6838 => "000000000000000000000000",
6839 => "000000000000000000000000",
6840 => "000000000000000000000000",
6841 => "000000000000000000000000",
6842 => "000000000000000000000000",
6843 => "000000000000000000000000",
6844 => "000000000000000000000000",
6845 => "000000000000000000000000",
6846 => "000000000000000000000000",
6847 => "000000000000000000000000",
6848 => "000000000000000000000000",
6849 => "000000000000000000000000",
6850 => "000000000000000000000000",
6851 => "000000000000000000000000",
6852 => "000000000000000000000000",
6853 => "000000000000000000000000",
6854 => "000000000000000000000000",
6855 => "000000000000000000000000",
6856 => "000000000000000000000000",
6857 => "000000000000000000000000",
6858 => "000000000000000000000000",
6859 => "000000000000000000000000",
6860 => "000000000000000000000000",
6861 => "000000000000000000000000",
6862 => "000000000000000000000000",
6863 => "000000000000000000000000",
6864 => "000000000000000000000000",
6865 => "000000000000000000000000",
6866 => "000000000000000000000000",
6867 => "000000000000000000000000",
6868 => "000000000000000000000000",
6869 => "000000000000000000000000",
6870 => "000000000000000000000000",
6871 => "000000000000000000000000",
6872 => "000000000000000000000000",
6873 => "000000000000000000000000",
6874 => "000000000000000000000000",
6875 => "000000000000000000000000",
6876 => "000000000000000000000000",
6877 => "000000000000000000000000",
6878 => "000000000000000000000000",
6879 => "000000000000000000000000",
6880 => "000000000000000000000000",
6881 => "000000000000000000000000",
6882 => "000000000000000000000000",
6883 => "000000000000000000000000",
6884 => "000000000000000000000000",
6885 => "000000000000000000000000",
6886 => "000000000000000000000000",
6887 => "000000000000000000000000",
6888 => "000000000000000000000000",
6889 => "000000000000000000000000",
6890 => "000000000000000000000000",
6891 => "000000000000000000000000",
6892 => "000000000000000000000000",
6893 => "000000000000000000000000",
6894 => "000000000000000000000000",
6895 => "000000000000000000000000",
6896 => "000000000000000000000000",
6897 => "000000000000000000000000",
6898 => "000000000000000000000000",
6899 => "000000000000000000000000",
6900 => "000000000000000000000000",
6901 => "000000000000000000000000",
6902 => "000000000000000000000000",
6903 => "000000000000000000000000",
6904 => "000000000000000000000000",
6905 => "000000000000000000000000",
6906 => "000000000000000000000000",
6907 => "000000000000000000000000",
6908 => "000000000000000000000000",
6909 => "000000000000000000000000",
6910 => "000000000000000000000000",
6911 => "000000000000000000000000",
6912 => "000000000000000000000000",
6913 => "000000000000000000000000",
6914 => "000000000000000000000000",
6915 => "000000000000000000000000",
6916 => "000000000000000000000000",
6917 => "000000000000000000000000",
6918 => "000000000000000000000000",
6919 => "000000000000000000000000",
6920 => "000000000000000000000000",
6921 => "000000000000000000000000",
6922 => "000000000000000000000000",
6923 => "000000000000000000000000",
6924 => "000000000000000000000000",
6925 => "000000000000000000000000",
6926 => "000000000000000000000000",
6927 => "000000000000000000000000",
6928 => "000000000000000000000000",
6929 => "000000000000000000000000",
6930 => "000000000000000000000000",
6931 => "000000000000000000000000",
6932 => "000000000000000000000000",
6933 => "000000000000000000000000",
6934 => "000000000000000000000000",
6935 => "000000000000000000000000",
6936 => "000000000000000000000000",
6937 => "000000000000000000000000",
6938 => "000000000000000000000000",
6939 => "000000000000000000000000",
6940 => "000000000000000000000000",
6941 => "000000000000000000000000",
6942 => "000000000000000000000000",
6943 => "000000000000000000000000",
6944 => "000000000000000000000000",
6945 => "000000000000000000000000",
6946 => "000000000000000000000000",
6947 => "000000000000000000000000",
6948 => "000000000000000000000000",
6949 => "000000000000000000000000",
6950 => "000000000000000000000000",
6951 => "000000000000000000000000",
6952 => "000000000000000000000000",
6953 => "000000000000000000000000",
6954 => "000000000000000000000000",
6955 => "000000000000000000000000",
6956 => "000000000000000000000000",
6957 => "000000000000000000000000",
6958 => "000000000000000000000000",
6959 => "000000000000000000000000",
6960 => "000001000000010000000100",
6961 => "010000110100001101000011",
6962 => "010000110100001101000011",
6963 => "000100100001001000010010",
6964 => "000000000000000000000000",
6965 => "001101000100000101001100",
6966 => "100010111010110011001011",
6967 => "100010111010110011001011",
6968 => "100010111010110011001011",
6969 => "100010111010110011001011",
6970 => "100010111010110011001011",
6971 => "100010111010110011001011",
6972 => "010110110111000110000101",
6973 => "000000000000000000000000",
6974 => "000000000000000000000000",
6975 => "010000110100001101000011",
6976 => "010000110100001101000011",
6977 => "000101110001011100010111",
6978 => "000000000000000000000000",
6979 => "000000000000000000000000",
6980 => "000000000000000000000000",
6981 => "000000000000000000000000",
6982 => "000000000000000000000000",
6983 => "000000000000000000000000",
6984 => "000000000000000000000000",
6985 => "000000000000000000000000",
6986 => "000000000000000000000000",
6987 => "000000000000000000000000",
6988 => "000000000000000000000000",
6989 => "000000000000000000000000",
6990 => "000000000000000000000000",
6991 => "000000000000000000000000",
6992 => "000000000000000000000000",
6993 => "000000000000000000000000",
6994 => "000000000000000000000000",
6995 => "000000000000000000000000",
6996 => "000000000000000000000000",
6997 => "000000000000000000000000",
6998 => "000000000000000000000000",
6999 => "000000000000000000000000",
7000 => "000000000000000000000000",
7001 => "000000000000000000000000",
7002 => "000000000000000000000000",
7003 => "000000000000000000000000",
7004 => "000000000000000000000000",
7005 => "000000000000000000000000",
7006 => "000000000000000000000000",
7007 => "000000000000000000000000",
7008 => "000000000000000000000000",
7009 => "000000000000000000000000",
7010 => "000000000000000000000000",
7011 => "000000000000000000000000",
7012 => "000000000000000000000000",
7013 => "000000000000000000000000",
7014 => "000000000000000000000000",
7015 => "000000000000000000000000",
7016 => "000000000000000000000000",
7017 => "000000000000000000000000",
7018 => "000000000000000000000000",
7019 => "000000000000000000000000",
7020 => "000000000000000000000000",
7021 => "000000000000000000000000",
7022 => "000000000000000000000000",
7023 => "000000000000000000000000",
7024 => "000000000000000000000000",
7025 => "000000000000000000000000",
7026 => "000000000000000000000000",
7027 => "000000000000000000000000",
7028 => "000000000000000000000000",
7029 => "000000000000000000000000",
7030 => "000000000000000000000000",
7031 => "000000000000000000000000",
7032 => "000000000000000000000000",
7033 => "000000000000000000000000",
7034 => "000000000000000000000000",
7035 => "000000000000000000000000",
7036 => "000000000000000000000000",
7037 => "000000000000000000000000",
7038 => "000000000000000000000000",
7039 => "000000000000000000000000",
7040 => "000000000000000000000000",
7041 => "000000000000000000000000",
7042 => "000000000000000000000000",
7043 => "000000000000000000000000",
7044 => "000000000000000000000000",
7045 => "000000000000000000000000",
7046 => "000000000000000000000000",
7047 => "000000000000000000000000",
7048 => "000000000000000000000000",
7049 => "000000000000000000000000",
7050 => "000000000000000000000000",
7051 => "000000000000000000000000",
7052 => "000000000000000000000000",
7053 => "000000000000000000000000",
7054 => "000000000000000000000000",
7055 => "000000000000000000000000",
7056 => "000000000000000000000000",
7057 => "000000000000000000000000",
7058 => "000000000000000000000000",
7059 => "000000000000000000000000",
7060 => "000000000000000000000000",
7061 => "000000000000000000000000",
7062 => "000000000000000000000000",
7063 => "000000000000000000000000",
7064 => "000000000000000000000000",
7065 => "000000000000000000000000",
7066 => "000000000000000000000000",
7067 => "000000000000000000000000",
7068 => "000000000000000000000000",
7069 => "000000000000000000000000",
7070 => "000000000000000000000000",
7071 => "000000000000000000000000",
7072 => "000000000000000000000000",
7073 => "000000000000000000000000",
7074 => "000000000000000000000000",
7075 => "000000000000000000000000",
7076 => "000000000000000000000000",
7077 => "000000000000000000000000",
7078 => "000000000000000000000000",
7079 => "000000000000000000000000",
7080 => "000000000000000000000000",
7081 => "000000000000000000000000",
7082 => "000000000000000000000000",
7083 => "000000000000000000000000",
7084 => "000000000000000000000000",
7085 => "000000000000000000000000",
7086 => "000000000000000000000000",
7087 => "000000000000000000000000",
7088 => "000000000000000000000000",
7089 => "000000000000000000000000",
7090 => "000000000000000000000000",
7091 => "000000000000000000000000",
7092 => "000000000000000000000000",
7093 => "000000000000000000000000",
7094 => "000000000000000000000000",
7095 => "000000000000000000000000",
7096 => "000000000000000000000000",
7097 => "000000000000000000000000",
7098 => "000000000000000000000000",
7099 => "000000000000000000000000",
7100 => "000000000000000000000000",
7101 => "000000000000000000000000",
7102 => "000000000000000000000000",
7103 => "000000000000000000000000",
7104 => "000000000000000000000000",
7105 => "000000000000000000000000",
7106 => "000000000000000000000000",
7107 => "000000000000000000000000",
7108 => "000000000000000000000000",
7109 => "000000000000000000000000",
7110 => "000001000000010000000100",
7111 => "010000110100001101000011",
7112 => "010000110100001101000011",
7113 => "000100100001001000010010",
7114 => "000000000000000000000000",
7115 => "000000000000000000000000",
7116 => "000000000000000000000000",
7117 => "000000000000000000000000",
7118 => "000000000000000000000000",
7119 => "000000000000000000000000",
7120 => "000000000000000000000000",
7121 => "000000000000000000000000",
7122 => "000000000000000000000000",
7123 => "000000000000000000000000",
7124 => "000000000000000000000000",
7125 => "010000110100001101000011",
7126 => "010000110100001101000011",
7127 => "000101110001011100010111",
7128 => "000000000000000000000000",
7129 => "000000000000000000000000",
7130 => "000000000000000000000000",
7131 => "000000000000000000000000",
7132 => "000000000000000000000000",
7133 => "000000000000000000000000",
7134 => "000000000000000000000000",
7135 => "000000000000000000000000",
7136 => "000000000000000000000000",
7137 => "000000000000000000000000",
7138 => "000000000000000000000000",
7139 => "000000000000000000000000",
7140 => "000000000000000000000000",
7141 => "000000000000000000000000",
7142 => "000000000000000000000000",
7143 => "000000000000000000000000",
7144 => "000000000000000000000000",
7145 => "000000000000000000000000",
7146 => "000000000000000000000000",
7147 => "000000000000000000000000",
7148 => "000000000000000000000000",
7149 => "000000000000000000000000",
7150 => "000000000000000000000000",
7151 => "000000000000000000000000",
7152 => "000000000000000000000000",
7153 => "000000000000000000000000",
7154 => "000000000000000000000000",
7155 => "000000000000000000000000",
7156 => "000000000000000000000000",
7157 => "000000000000000000000000",
7158 => "000000000000000000000000",
7159 => "000000000000000000000000",
7160 => "000000000000000000000000",
7161 => "000000000000000000000000",
7162 => "000000000000000000000000",
7163 => "000000000000000000000000",
7164 => "000000000000000000000000",
7165 => "000000000000000000000000",
7166 => "000000000000000000000000",
7167 => "000000000000000000000000",
7168 => "000000000000000000000000",
7169 => "000000000000000000000000",
7170 => "000000000000000000000000",
7171 => "000000000000000000000000",
7172 => "000000000000000000000000",
7173 => "000000000000000000000000",
7174 => "000000000000000000000000",
7175 => "000000000000000000000000",
7176 => "000000000000000000000000",
7177 => "000000000000000000000000",
7178 => "000000000000000000000000",
7179 => "000000000000000000000000",
7180 => "000000000000000000000000",
7181 => "000000000000000000000000",
7182 => "000000000000000000000000",
7183 => "000000000000000000000000",
7184 => "000000000000000000000000",
7185 => "000000000000000000000000",
7186 => "000000000000000000000000",
7187 => "000000000000000000000000",
7188 => "000000000000000000000000",
7189 => "000000000000000000000000",
7190 => "000000000000000000000000",
7191 => "000000000000000000000000",
7192 => "000000000000000000000000",
7193 => "000000000000000000000000",
7194 => "000000000000000000000000",
7195 => "000000000000000000000000",
7196 => "000000000000000000000000",
7197 => "000000000000000000000000",
7198 => "000000000000000000000000",
7199 => "000000000000000000000000",
7200 => "000000000000000000000000",
7201 => "000000000000000000000000",
7202 => "000000000000000000000000",
7203 => "000000000000000000000000",
7204 => "000000000000000000000000",
7205 => "000000000000000000000000",
7206 => "000000000000000000000000",
7207 => "000000000000000000000000",
7208 => "000000000000000000000000",
7209 => "000000000000000000000000",
7210 => "000000000000000000000000",
7211 => "000000000000000000000000",
7212 => "000000000000000000000000",
7213 => "000000000000000000000000",
7214 => "000000000000000000000000",
7215 => "000000000000000000000000",
7216 => "000000000000000000000000",
7217 => "000000000000000000000000",
7218 => "000000000000000000000000",
7219 => "000000000000000000000000",
7220 => "000000000000000000000000",
7221 => "000000000000000000000000",
7222 => "000000000000000000000000",
7223 => "000000000000000000000000",
7224 => "000000000000000000000000",
7225 => "000000000000000000000000",
7226 => "000000000000000000000000",
7227 => "000000000000000000000000",
7228 => "000000000000000000000000",
7229 => "000000000000000000000000",
7230 => "000000000000000000000000",
7231 => "000000000000000000000000",
7232 => "000000000000000000000000",
7233 => "000000000000000000000000",
7234 => "000000000000000000000000",
7235 => "000000000000000000000000",
7236 => "000000000000000000000000",
7237 => "000000000000000000000000",
7238 => "000000000000000000000000",
7239 => "000000000000000000000000",
7240 => "000000000000000000000000",
7241 => "000000000000000000000000",
7242 => "000000000000000000000000",
7243 => "000000000000000000000000",
7244 => "000000000000000000000000",
7245 => "000000000000000000000000",
7246 => "000000000000000000000000",
7247 => "000000000000000000000000",
7248 => "000000000000000000000000",
7249 => "000000000000000000000000",
7250 => "000000000000000000000000",
7251 => "000000000000000000000000",
7252 => "000000000000000000000000",
7253 => "000000000000000000000000",
7254 => "000000000000000000000000",
7255 => "000000000000000000000000",
7256 => "000000000000000000000000",
7257 => "000000000000000000000000",
7258 => "000000000000000000000000",
7259 => "000000000000000000000000",
7260 => "000001000000010000000100",
7261 => "010000110100001101000011",
7262 => "010000110100001101000011",
7263 => "000100100001001000010010",
7264 => "000000000000000000000000",
7265 => "000000000000000000000000",
7266 => "000000000000000000000000",
7267 => "000000000000000000000000",
7268 => "000000000000000000000000",
7269 => "000000000000000000000000",
7270 => "000000000000000000000000",
7271 => "000000000000000000000000",
7272 => "000000000000000000000000",
7273 => "000000000000000000000000",
7274 => "000000000000000000000000",
7275 => "010000110100001101000011",
7276 => "010000110100001101000011",
7277 => "000101110001011100010111",
7278 => "000000000000000000000000",
7279 => "000000000000000000000000",
7280 => "000000000000000000000000",
7281 => "000000000000000000000000",
7282 => "000000000000000000000000",
7283 => "000000000000000000000000",
7284 => "000000000000000000000000",
7285 => "000000000000000000000000",
7286 => "000000000000000000000000",
7287 => "000000000000000000000000",
7288 => "000000000000000000000000",
7289 => "000000000000000000000000",
7290 => "000000000000000000000000",
7291 => "000000000000000000000000",
7292 => "000000000000000000000000",
7293 => "000000000000000000000000",
7294 => "000000000000000000000000",
7295 => "000000000000000000000000",
7296 => "000000000000000000000000",
7297 => "000000000000000000000000",
7298 => "000000000000000000000000",
7299 => "000000000000000000000000",
7300 => "000000000000000000000000",
7301 => "000000000000000000000000",
7302 => "000000000000000000000000",
7303 => "000000000000000000000000",
7304 => "000000000000000000000000",
7305 => "000000000000000000000000",
7306 => "000000000000000000000000",
7307 => "000000000000000000000000",
7308 => "000000000000000000000000",
7309 => "000000000000000000000000",
7310 => "000000000000000000000000",
7311 => "000000000000000000000000",
7312 => "000000000000000000000000",
7313 => "000000000000000000000000",
7314 => "000000000000000000000000",
7315 => "000000000000000000000000",
7316 => "000000000000000000000000",
7317 => "000000000000000000000000",
7318 => "000000000000000000000000",
7319 => "000000000000000000000000",
7320 => "000000000000000000000000",
7321 => "000000000000000000000000",
7322 => "000000000000000000000000",
7323 => "000000000000000000000000",
7324 => "000000000000000000000000",
7325 => "000000000000000000000000",
7326 => "000000000000000000000000",
7327 => "000000000000000000000000",
7328 => "000000000000000000000000",
7329 => "000000000000000000000000",
7330 => "000000000000000000000000",
7331 => "000000000000000000000000",
7332 => "000000000000000000000000",
7333 => "000000000000000000000000",
7334 => "000000000000000000000000",
7335 => "000000000000000000000000",
7336 => "000000000000000000000000",
7337 => "000000000000000000000000",
7338 => "000000000000000000000000",
7339 => "000000000000000000000000",
7340 => "000000000000000000000000",
7341 => "000000000000000000000000",
7342 => "000000000000000000000000",
7343 => "000000000000000000000000",
7344 => "000000000000000000000000",
7345 => "000000000000000000000000",
7346 => "000000000000000000000000",
7347 => "000000000000000000000000",
7348 => "000000000000000000000000",
7349 => "000000000000000000000000",
7350 => "000000000000000000000000",
7351 => "000000000000000000000000",
7352 => "000000000000000000000000",
7353 => "000000000000000000000000",
7354 => "000000000000000000000000",
7355 => "000000000000000000000000",
7356 => "000000000000000000000000",
7357 => "000000000000000000000000",
7358 => "000000000000000000000000",
7359 => "000000000000000000000000",
7360 => "000000000000000000000000",
7361 => "000000000000000000000000",
7362 => "000000000000000000000000",
7363 => "000000000000000000000000",
7364 => "000000000000000000000000",
7365 => "000000000000000000000000",
7366 => "000000000000000000000000",
7367 => "000000000000000000000000",
7368 => "000000000000000000000000",
7369 => "000000000000000000000000",
7370 => "000000000000000000000000",
7371 => "000000000000000000000000",
7372 => "000000000000000000000000",
7373 => "000000000000000000000000",
7374 => "000000000000000000000000",
7375 => "000000000000000000000000",
7376 => "000000000000000000000000",
7377 => "000000000000000000000000",
7378 => "000000000000000000000000",
7379 => "000000000000000000000000",
7380 => "000000000000000000000000",
7381 => "000000000000000000000000",
7382 => "000000000000000000000000",
7383 => "000000000000000000000000",
7384 => "000000000000000000000000",
7385 => "000000000000000000000000",
7386 => "000000000000000000000000",
7387 => "000000000000000000000000",
7388 => "000000000000000000000000",
7389 => "000000000000000000000000",
7390 => "000000000000000000000000",
7391 => "000000000000000000000000",
7392 => "000000000000000000000000",
7393 => "000000000000000000000000",
7394 => "000000000000000000000000",
7395 => "000000000000000000000000",
7396 => "000000000000000000000000",
7397 => "000000000000000000000000",
7398 => "000000000000000000000000",
7399 => "000000000000000000000000",
7400 => "000000000000000000000000",
7401 => "000000000000000000000000",
7402 => "000000000000000000000000",
7403 => "000000000000000000000000",
7404 => "000000000000000000000000",
7405 => "000000000000000000000000",
7406 => "000000000000000000000000",
7407 => "000000000000000000000000",
7408 => "000000000000000000000000",
7409 => "000000000000000000000000",
7410 => "000001000000010000000100",
7411 => "010000110100001101000011",
7412 => "010000110100001101000011",
7413 => "000100100001001000010010",
7414 => "000000000000000000000000",
7415 => "001100100011111001001001",
7416 => "100001011010010111000010",
7417 => "100001011010010111000010",
7418 => "100001011010010111000010",
7419 => "100001011010010111000010",
7420 => "100001011010010111000010",
7421 => "100001011010010111000010",
7422 => "010101110110110001111111",
7423 => "000000000000000000000000",
7424 => "000000000000000000000000",
7425 => "010000110100001101000011",
7426 => "010000110100001101000011",
7427 => "000101110001011100010111",
7428 => "000000000000000000000000",
7429 => "000000000000000000000000",
7430 => "000000000000000000000000",
7431 => "000000000000000000000000",
7432 => "000000000000000000000000",
7433 => "000000000000000000000000",
7434 => "000000000000000000000000",
7435 => "000000000000000000000000",
7436 => "000000000000000000000000",
7437 => "000000000000000000000000",
7438 => "000000000000000000000000",
7439 => "000000000000000000000000",
7440 => "000000000000000000000000",
7441 => "000000000000000000000000",
7442 => "000000000000000000000000",
7443 => "000000000000000000000000",
7444 => "000000000000000000000000",
7445 => "000000000000000000000000",
7446 => "000000000000000000000000",
7447 => "000000000000000000000000",
7448 => "000000000000000000000000",
7449 => "000000000000000000000000",
7450 => "000000000000000000000000",
7451 => "000000000000000000000000",
7452 => "000000000000000000000000",
7453 => "000000000000000000000000",
7454 => "000000000000000000000000",
7455 => "000000000000000000000000",
7456 => "000000000000000000000000",
7457 => "000000000000000000000000",
7458 => "000000000000000000000000",
7459 => "000000000000000000000000",
7460 => "000000000000000000000000",
7461 => "000000000000000000000000",
7462 => "000000000000000000000000",
7463 => "000000000000000000000000",
7464 => "000000000000000000000000",
7465 => "000000000000000000000000",
7466 => "000000000000000000000000",
7467 => "000000000000000000000000",
7468 => "000000000000000000000000",
7469 => "000000000000000000000000",
7470 => "000000000000000000000000",
7471 => "000000000000000000000000",
7472 => "000000000000000000000000",
7473 => "000000000000000000000000",
7474 => "000000000000000000000000",
7475 => "000000000000000000000000",
7476 => "000000000000000000000000",
7477 => "000000000000000000000000",
7478 => "000000000000000000000000",
7479 => "000000000000000000000000",
7480 => "000000000000000000000000",
7481 => "000000000000000000000000",
7482 => "000000000000000000000000",
7483 => "000000000000000000000000",
7484 => "000000000000000000000000",
7485 => "000000000000000000000000",
7486 => "000000000000000000000000",
7487 => "000000000000000000000000",
7488 => "000000000000000000000000",
7489 => "000000000000000000000000",
7490 => "000000000000000000000000",
7491 => "000000000000000000000000",
7492 => "000000000000000000000000",
7493 => "000000000000000000000000",
7494 => "000000000000000000000000",
7495 => "000000000000000000000000",
7496 => "000000000000000000000000",
7497 => "000000000000000000000000",
7498 => "000000000000000000000000",
7499 => "000000000000000000000000",
7500 => "000000000000000000000000",
7501 => "000000000000000000000000",
7502 => "000000000000000000000000",
7503 => "000000000000000000000000",
7504 => "000000000000000000000000",
7505 => "000000000000000000000000",
7506 => "000000000000000000000000",
7507 => "000000000000000000000000",
7508 => "000000000000000000000000",
7509 => "000000000000000000000000",
7510 => "000000000000000000000000",
7511 => "000000000000000000000000",
7512 => "000000000000000000000000",
7513 => "000000000000000000000000",
7514 => "000000000000000000000000",
7515 => "000000000000000000000000",
7516 => "000000000000000000000000",
7517 => "000000000000000000000000",
7518 => "000000000000000000000000",
7519 => "000000000000000000000000",
7520 => "000000000000000000000000",
7521 => "000000000000000000000000",
7522 => "000000000000000000000000",
7523 => "000000000000000000000000",
7524 => "000000000000000000000000",
7525 => "000000000000000000000000",
7526 => "000000000000000000000000",
7527 => "000000000000000000000000",
7528 => "000000000000000000000000",
7529 => "000000000000000000000000",
7530 => "000000000000000000000000",
7531 => "000000000000000000000000",
7532 => "000000000000000000000000",
7533 => "000000000000000000000000",
7534 => "000000000000000000000000",
7535 => "000000000000000000000000",
7536 => "000000000000000000000000",
7537 => "000000000000000000000000",
7538 => "000000000000000000000000",
7539 => "000000000000000000000000",
7540 => "000000000000000000000000",
7541 => "000000000000000000000000",
7542 => "000000000000000000000000",
7543 => "000000000000000000000000",
7544 => "000000000000000000000000",
7545 => "000000000000000000000000",
7546 => "000000000000000000000000",
7547 => "000000000000000000000000",
7548 => "000000000000000000000000",
7549 => "000000000000000000000000",
7550 => "000000000000000000000000",
7551 => "000000000000000000000000",
7552 => "000000000000000000000000",
7553 => "000000000000000000000000",
7554 => "000000000000000000000000",
7555 => "000000000000000000000000",
7556 => "000000000000000000000000",
7557 => "000000000000000000000000",
7558 => "000000000000000000000000",
7559 => "000000000000000000000000",
7560 => "000001000000010000000100",
7561 => "010000110100001101000011",
7562 => "010000110100001101000011",
7563 => "000100100001001000010010",
7564 => "000000000000000000000000",
7565 => "001111000100101001010111",
7566 => "100111111100010111101000",
7567 => "100111111100010111101000",
7568 => "100111111100010111101000",
7569 => "100111111100010111101000",
7570 => "100111111100010111101000",
7571 => "100111111100010111101000",
7572 => "011010001000000110011000",
7573 => "000000000000000000000000",
7574 => "000000000000000000000000",
7575 => "010000110100001101000011",
7576 => "010000110100001101000011",
7577 => "000101110001011100010111",
7578 => "000000000000000000000000",
7579 => "000000000000000000000000",
7580 => "000000000000000000000000",
7581 => "000000000000000000000000",
7582 => "000000000000000000000000",
7583 => "000000000000000000000000",
7584 => "000000000000000000000000",
7585 => "000000000000000000000000",
7586 => "000000000000000000000000",
7587 => "000000000000000000000000",
7588 => "000000000000000000000000",
7589 => "000000000000000000000000",
7590 => "000000000000000000000000",
7591 => "000000000000000000000000",
7592 => "000000000000000000000000",
7593 => "000000000000000000000000",
7594 => "000000000000000000000000",
7595 => "000000000000000000000000",
7596 => "000000000000000000000000",
7597 => "000000000000000000000000",
7598 => "000000000000000000000000",
7599 => "000000000000000000000000",
7600 => "000000000000000000000000",
7601 => "000000000000000000000000",
7602 => "000000000000000000000000",
7603 => "000000000000000000000000",
7604 => "000000000000000000000000",
7605 => "000000000000000000000000",
7606 => "000000000000000000000000",
7607 => "000000000000000000000000",
7608 => "000000000000000000000000",
7609 => "000000000000000000000000",
7610 => "000000000000000000000000",
7611 => "000000000000000000000000",
7612 => "000000000000000000000000",
7613 => "000000000000000000000000",
7614 => "000000000000000000000000",
7615 => "000000000000000000000000",
7616 => "000000000000000000000000",
7617 => "000000000000000000000000",
7618 => "000000000000000000000000",
7619 => "000000000000000000000000",
7620 => "000000000000000000000000",
7621 => "000000000000000000000000",
7622 => "000000000000000000000000",
7623 => "000000000000000000000000",
7624 => "000000000000000000000000",
7625 => "000000000000000000000000",
7626 => "000000000000000000000000",
7627 => "000000000000000000000000",
7628 => "000000000000000000000000",
7629 => "000000000000000000000000",
7630 => "000000000000000000000000",
7631 => "000000000000000000000000",
7632 => "000000000000000000000000",
7633 => "000000000000000000000000",
7634 => "000000000000000000000000",
7635 => "000000000000000000000000",
7636 => "000000000000000000000000",
7637 => "000000000000000000000000",
7638 => "000000000000000000000000",
7639 => "000000000000000000000000",
7640 => "000000000000000000000000",
7641 => "000000000000000000000000",
7642 => "000000000000000000000000",
7643 => "000000000000000000000000",
7644 => "000000000000000000000000",
7645 => "000000000000000000000000",
7646 => "000000000000000000000000",
7647 => "000000000000000000000000",
7648 => "000000000000000000000000",
7649 => "000000000000000000000000",
7650 => "000000000000000000000000",
7651 => "000000000000000000000000",
7652 => "000000000000000000000000",
7653 => "000000000000000000000000",
7654 => "000000000000000000000000",
7655 => "000000000000000000000000",
7656 => "000000000000000000000000",
7657 => "000000000000000000000000",
7658 => "000000000000000000000000",
7659 => "000000000000000000000000",
7660 => "000000000000000000000000",
7661 => "000000000000000000000000",
7662 => "000000000000000000000000",
7663 => "000000000000000000000000",
7664 => "000000000000000000000000",
7665 => "000000000000000000000000",
7666 => "000000000000000000000000",
7667 => "000000000000000000000000",
7668 => "000000000000000000000000",
7669 => "000000000000000000000000",
7670 => "000000000000000000000000",
7671 => "000000000000000000000000",
7672 => "000000000000000000000000",
7673 => "000000000000000000000000",
7674 => "000000000000000000000000",
7675 => "000000000000000000000000",
7676 => "000000000000000000000000",
7677 => "000000000000000000000000",
7678 => "000000000000000000000000",
7679 => "000000000000000000000000",
7680 => "000000000000000000000000",
7681 => "000000000000000000000000",
7682 => "000000000000000000000000",
7683 => "000000000000000000000000",
7684 => "000000000000000000000000",
7685 => "000000000000000000000000",
7686 => "000000000000000000000000",
7687 => "000000000000000000000000",
7688 => "000000000000000000000000",
7689 => "000000000000000000000000",
7690 => "000000000000000000000000",
7691 => "000000000000000000000000",
7692 => "000000000000000000000000",
7693 => "000000000000000000000000",
7694 => "000000000000000000000000",
7695 => "000000000000000000000000",
7696 => "000000000000000000000000",
7697 => "000000000000000000000000",
7698 => "000000000000000000000000",
7699 => "000000000000000000000000",
7700 => "000000000000000000000000",
7701 => "000000000000000000000000",
7702 => "000000000000000000000000",
7703 => "000000000000000000000000",
7704 => "000000000000000000000000",
7705 => "000000000000000000000000",
7706 => "000000000000000000000000",
7707 => "000000000000000000000000",
7708 => "000011000000110000001100",
7709 => "000111010001110100011101",
7710 => "001000000010000000100000",
7711 => "010000110100001101000011",
7712 => "010000110100001101000011",
7713 => "000100100001001000010010",
7714 => "000000000000000000000000",
7715 => "001111000100101001010111",
7716 => "100111111100010111101000",
7717 => "100111111100010111101000",
7718 => "100111111100010111101000",
7719 => "100111111100010111101000",
7720 => "100111111100010111101000",
7721 => "100111111100010111101000",
7722 => "011010001000000110011000",
7723 => "000000000000000000000000",
7724 => "000000000000000000000000",
7725 => "010000110100001101000011",
7726 => "010000110100001101000011",
7727 => "001010100010101000101010",
7728 => "000111010001110100011101",
7729 => "000101000001010000010100",
7730 => "000000000000000000000000",
7731 => "000000000000000000000000",
7732 => "000000000000000000000000",
7733 => "000000000000000000000000",
7734 => "000000000000000000000000",
7735 => "000000000000000000000000",
7736 => "000000000000000000000000",
7737 => "000000000000000000000000",
7738 => "000000000000000000000000",
7739 => "000000000000000000000000",
7740 => "000000000000000000000000",
7741 => "000000000000000000000000",
7742 => "000000000000000000000000",
7743 => "000000000000000000000000",
7744 => "000000000000000000000000",
7745 => "000000000000000000000000",
7746 => "000000000000000000000000",
7747 => "000000000000000000000000",
7748 => "000000000000000000000000",
7749 => "000000000000000000000000",
7750 => "000000000000000000000000",
7751 => "000000000000000000000000",
7752 => "000000000000000000000000",
7753 => "000000000000000000000000",
7754 => "000000000000000000000000",
7755 => "000000000000000000000000",
7756 => "000000000000000000000000",
7757 => "000000000000000000000000",
7758 => "000000000000000000000000",
7759 => "000000000000000000000000",
7760 => "000000000000000000000000",
7761 => "000000000000000000000000",
7762 => "000000000000000000000000",
7763 => "000000000000000000000000",
7764 => "000000000000000000000000",
7765 => "000000000000000000000000",
7766 => "000000000000000000000000",
7767 => "000000000000000000000000",
7768 => "000000000000000000000000",
7769 => "000000000000000000000000",
7770 => "000000000000000000000000",
7771 => "000000000000000000000000",
7772 => "000000000000000000000000",
7773 => "000000000000000000000000",
7774 => "000000000000000000000000",
7775 => "000000000000000000000000",
7776 => "000000000000000000000000",
7777 => "000000000000000000000000",
7778 => "000000000000000000000000",
7779 => "000000000000000000000000",
7780 => "000000000000000000000000",
7781 => "000000000000000000000000",
7782 => "000000000000000000000000",
7783 => "000000000000000000000000",
7784 => "000000000000000000000000",
7785 => "000000000000000000000000",
7786 => "000000000000000000000000",
7787 => "000000000000000000000000",
7788 => "000000000000000000000000",
7789 => "000000000000000000000000",
7790 => "000000000000000000000000",
7791 => "000000000000000000000000",
7792 => "000000000000000000000000",
7793 => "000000000000000000000000",
7794 => "000000000000000000000000",
7795 => "000000000000000000000000",
7796 => "000000000000000000000000",
7797 => "000000000000000000000000",
7798 => "000000000000000000000000",
7799 => "000000000000000000000000",
7800 => "000000000000000000000000",
7801 => "000000000000000000000000",
7802 => "000000000000000000000000",
7803 => "000000000000000000000000",
7804 => "000000000000000000000000",
7805 => "000000000000000000000000",
7806 => "000000000000000000000000",
7807 => "000000000000000000000000",
7808 => "000000000000000000000000",
7809 => "000000000000000000000000",
7810 => "000000000000000000000000",
7811 => "000000000000000000000000",
7812 => "000000000000000000000000",
7813 => "000000000000000000000000",
7814 => "000000000000000000000000",
7815 => "000000000000000000000000",
7816 => "000000000000000000000000",
7817 => "000000000000000000000000",
7818 => "000000000000000000000000",
7819 => "000000000000000000000000",
7820 => "000000000000000000000000",
7821 => "000000000000000000000000",
7822 => "000000000000000000000000",
7823 => "000000000000000000000000",
7824 => "000000000000000000000000",
7825 => "000000000000000000000000",
7826 => "000000000000000000000000",
7827 => "000000000000000000000000",
7828 => "000000000000000000000000",
7829 => "000000000000000000000000",
7830 => "000000000000000000000000",
7831 => "000000000000000000000000",
7832 => "000000000000000000000000",
7833 => "000000000000000000000000",
7834 => "000000000000000000000000",
7835 => "000000000000000000000000",
7836 => "000000000000000000000000",
7837 => "000000000000000000000000",
7838 => "000000000000000000000000",
7839 => "000000000000000000000000",
7840 => "000000000000000000000000",
7841 => "000000000000000000000000",
7842 => "000000000000000000000000",
7843 => "000000000000000000000000",
7844 => "000000000000000000000000",
7845 => "000000000000000000000000",
7846 => "000000000000000000000000",
7847 => "000000000000000000000000",
7848 => "000000000000000000000000",
7849 => "000000000000000000000000",
7850 => "000000000000000000000000",
7851 => "000000000000000000000000",
7852 => "000000000000000000000000",
7853 => "000000000000000000000000",
7854 => "000000000000000000000000",
7855 => "000000000000000000000000",
7856 => "000000000000000000000000",
7857 => "000000000000000000000000",
7858 => "000110110001101100011011",
7859 => "010000110100001101000011",
7860 => "010000110100001101000011",
7861 => "010000110100001101000011",
7862 => "010000110100001101000011",
7863 => "000100100001001000010010",
7864 => "000000000000000000000000",
7865 => "001111000100101001010111",
7866 => "100111111100010111101000",
7867 => "100111111100010111101000",
7868 => "100111111100010111101000",
7869 => "100111111100010111101000",
7870 => "100111111100010111101000",
7871 => "100111111100010111101000",
7872 => "011010001000000110011000",
7873 => "000000000000000000000000",
7874 => "000000000000000000000000",
7875 => "010000110100001101000011",
7876 => "010000110100001101000011",
7877 => "010000110100001101000011",
7878 => "010000110100001101000011",
7879 => "001011100010111000101110",
7880 => "000000000000000000000000",
7881 => "000000000000000000000000",
7882 => "000000000000000000000000",
7883 => "000000000000000000000000",
7884 => "000000000000000000000000",
7885 => "000000000000000000000000",
7886 => "000000000000000000000000",
7887 => "000000000000000000000000",
7888 => "000000000000000000000000",
7889 => "000000000000000000000000",
7890 => "000000000000000000000000",
7891 => "000000000000000000000000",
7892 => "000000000000000000000000",
7893 => "000000000000000000000000",
7894 => "000000000000000000000000",
7895 => "000000000000000000000000",
7896 => "000000000000000000000000",
7897 => "000000000000000000000000",
7898 => "000000000000000000000000",
7899 => "000000000000000000000000",
7900 => "000000000000000000000000",
7901 => "000000000000000000000000",
7902 => "000000000000000000000000",
7903 => "000000000000000000000000",
7904 => "000000000000000000000000",
7905 => "000000000000000000000000",
7906 => "000000000000000000000000",
7907 => "000000000000000000000000",
7908 => "000000000000000000000000",
7909 => "000000000000000000000000",
7910 => "000000000000000000000000",
7911 => "000000000000000000000000",
7912 => "000000000000000000000000",
7913 => "000000000000000000000000",
7914 => "000000000000000000000000",
7915 => "000000000000000000000000",
7916 => "000000000000000000000000",
7917 => "000000000000000000000000",
7918 => "000000000000000000000000",
7919 => "000000000000000000000000",
7920 => "000000000000000000000000",
7921 => "000000000000000000000000",
7922 => "000000000000000000000000",
7923 => "000000000000000000000000",
7924 => "000000000000000000000000",
7925 => "000000000000000000000000",
7926 => "000000000000000000000000",
7927 => "000000000000000000000000",
7928 => "000000000000000000000000",
7929 => "000000000000000000000000",
7930 => "000000000000000000000000",
7931 => "000000000000000000000000",
7932 => "000000000000000000000000",
7933 => "000000000000000000000000",
7934 => "000000000000000000000000",
7935 => "000000000000000000000000",
7936 => "000000000000000000000000",
7937 => "000000000000000000000000",
7938 => "000000000000000000000000",
7939 => "000000000000000000000000",
7940 => "000000000000000000000000",
7941 => "000000000000000000000000",
7942 => "000000000000000000000000",
7943 => "000000000000000000000000",
7944 => "000000000000000000000000",
7945 => "000000000000000000000000",
7946 => "000000000000000000000000",
7947 => "000000000000000000000000",
7948 => "000000000000000000000000",
7949 => "000000000000000000000000",
7950 => "000000000000000000000000",
7951 => "000000000000000000000000",
7952 => "000000000000000000000000",
7953 => "000000000000000000000000",
7954 => "000000000000000000000000",
7955 => "000000000000000000000000",
7956 => "000000000000000000000000",
7957 => "000000000000000000000000",
7958 => "000000000000000000000000",
7959 => "000000000000000000000000",
7960 => "000000000000000000000000",
7961 => "000000000000000000000000",
7962 => "000000000000000000000000",
7963 => "000000000000000000000000",
7964 => "000000000000000000000000",
7965 => "000000000000000000000000",
7966 => "000000000000000000000000",
7967 => "000000000000000000000000",
7968 => "000000000000000000000000",
7969 => "000000000000000000000000",
7970 => "000000000000000000000000",
7971 => "000000000000000000000000",
7972 => "000000000000000000000000",
7973 => "000000000000000000000000",
7974 => "000000000000000000000000",
7975 => "000000000000000000000000",
7976 => "000000000000000000000000",
7977 => "000000000000000000000000",
7978 => "000000000000000000000000",
7979 => "000000000000000000000000",
7980 => "000000000000000000000000",
7981 => "000000000000000000000000",
7982 => "000000000000000000000000",
7983 => "000000000000000000000000",
7984 => "000000000000000000000000",
7985 => "000000000000000000000000",
7986 => "000000000000000000000000",
7987 => "000000000000000000000000",
7988 => "000000000000000000000000",
7989 => "000000000000000000000000",
7990 => "000000000000000000000000",
7991 => "000000000000000000000000",
7992 => "000000000000000000000000",
7993 => "000000000000000000000000",
7994 => "000000000000000000000000",
7995 => "000000000000000000000000",
7996 => "000000000000000000000000",
7997 => "000000000000000000000000",
7998 => "000000000000000000000000",
7999 => "000000000000000000000000",
8000 => "000000000000000000000000",
8001 => "000000000000000000000000",
8002 => "000000000000000000000000",
8003 => "000000010000000100000001",
8004 => "000001100000011000000110",
8005 => "000001100000011000000110",
8006 => "000010010000100100001001",
8007 => "000010100000101000001010",
8008 => "000111100001111000011110",
8009 => "001111010011110100111101",
8010 => "001111010011110100111101",
8011 => "010000110100001101000011",
8012 => "010000110100001101000011",
8013 => "000100100001001000010010",
8014 => "000000000000000000000000",
8015 => "001111000100101001010111",
8016 => "100111111100010111101000",
8017 => "100111111100010111101000",
8018 => "100111111100010111101000",
8019 => "100111111100010111101000",
8020 => "100111111100010111101000",
8021 => "100111111100010111101000",
8022 => "011010001000000110011000",
8023 => "000000000000000000000000",
8024 => "000000000000000000000000",
8025 => "010000110100001101000011",
8026 => "010000110100001101000011",
8027 => "001111110011111100111111",
8028 => "001111010011110100111101",
8029 => "001011010010110100101101",
8030 => "000010100000101000001010",
8031 => "000010100000101000001010",
8032 => "000001100000011000000110",
8033 => "000001100000011000000110",
8034 => "000000100000001000000010",
8035 => "000000000000000000000000",
8036 => "000000000000000000000000",
8037 => "000000000000000000000000",
8038 => "000000000000000000000000",
8039 => "000000000000000000000000",
8040 => "000000000000000000000000",
8041 => "000000000000000000000000",
8042 => "000000000000000000000000",
8043 => "000000000000000000000000",
8044 => "000000000000000000000000",
8045 => "000000000000000000000000",
8046 => "000000000000000000000000",
8047 => "000000000000000000000000",
8048 => "000000000000000000000000",
8049 => "000000000000000000000000",
8050 => "000000000000000000000000",
8051 => "000000000000000000000000",
8052 => "000000000000000000000000",
8053 => "000000000000000000000000",
8054 => "000000000000000000000000",
8055 => "000000000000000000000000",
8056 => "000000000000000000000000",
8057 => "000000000000000000000000",
8058 => "000000000000000000000000",
8059 => "000000000000000000000000",
8060 => "000000000000000000000000",
8061 => "000000000000000000000000",
8062 => "000000000000000000000000",
8063 => "000000000000000000000000",
8064 => "000000000000000000000000",
8065 => "000000000000000000000000",
8066 => "000000000000000000000000",
8067 => "000000000000000000000000",
8068 => "000000000000000000000000",
8069 => "000000000000000000000000",
8070 => "000000000000000000000000",
8071 => "000000000000000000000000",
8072 => "000000000000000000000000",
8073 => "000000000000000000000000",
8074 => "000000000000000000000000",
8075 => "000000000000000000000000",
8076 => "000000000000000000000000",
8077 => "000000000000000000000000",
8078 => "000000000000000000000000",
8079 => "000000000000000000000000",
8080 => "000000000000000000000000",
8081 => "000000000000000000000000",
8082 => "000000000000000000000000",
8083 => "000000000000000000000000",
8084 => "000000000000000000000000",
8085 => "000000000000000000000000",
8086 => "000000000000000000000000",
8087 => "000000000000000000000000",
8088 => "000000000000000000000000",
8089 => "000000000000000000000000",
8090 => "000000000000000000000000",
8091 => "000000000000000000000000",
8092 => "000000000000000000000000",
8093 => "000000000000000000000000",
8094 => "000000000000000000000000",
8095 => "000000000000000000000000",
8096 => "000000000000000000000000",
8097 => "000000000000000000000000",
8098 => "000000000000000000000000",
8099 => "000000000000000000000000",
8100 => "000000000000000000000000",
8101 => "000000000000000000000000",
8102 => "000000000000000000000000",
8103 => "000000000000000000000000",
8104 => "000000000000000000000000",
8105 => "000000000000000000000000",
8106 => "000000000000000000000000",
8107 => "000000000000000000000000",
8108 => "000000000000000000000000",
8109 => "000000000000000000000000",
8110 => "000000000000000000000000",
8111 => "000000000000000000000000",
8112 => "000000000000000000000000",
8113 => "000000000000000000000000",
8114 => "000000000000000000000000",
8115 => "000000000000000000000000",
8116 => "000000000000000000000000",
8117 => "000000000000000000000000",
8118 => "000000000000000000000000",
8119 => "000000000000000000000000",
8120 => "000000000000000000000000",
8121 => "000000000000000000000000",
8122 => "000000000000000000000000",
8123 => "000000000000000000000000",
8124 => "000000000000000000000000",
8125 => "000000000000000000000000",
8126 => "000000000000000000000000",
8127 => "000000000000000000000000",
8128 => "000000000000000000000000",
8129 => "000000000000000000000000",
8130 => "000000000000000000000000",
8131 => "000000000000000000000000",
8132 => "000000000000000000000000",
8133 => "000000000000000000000000",
8134 => "000000000000000000000000",
8135 => "000000000000000000000000",
8136 => "000000000000000000000000",
8137 => "000000000000000000000000",
8138 => "000000000000000000000000",
8139 => "000000000000000000000000",
8140 => "000000000000000000000000",
8141 => "000000000000000000000000",
8142 => "000000000000000000000000",
8143 => "000000000000000000000000",
8144 => "000000000000000000000000",
8145 => "000000000000000000000000",
8146 => "000000000000000000000000",
8147 => "000000000000000000000000",
8148 => "000000000000000000000000",
8149 => "000000000000000000000000",
8150 => "000000000000000000000000",
8151 => "000000000000000000000000",
8152 => "000000000000000000000000",
8153 => "000001100000011000000110",
8154 => "010000110100001101000011",
8155 => "010000110100001101000011",
8156 => "010111110101111101011111",
8157 => "011001100110011001100110",
8158 => "001111010011110100111101",
8159 => "000000000000000000000000",
8160 => "000001000000010000000100",
8161 => "010000110100001101000011",
8162 => "010000110100001101000011",
8163 => "000100100001001000010010",
8164 => "000000000000000000000000",
8165 => "001111000100101001010111",
8166 => "100111111100010111101000",
8167 => "100111111100010111101000",
8168 => "100111111100010111101000",
8169 => "100111111100010111101000",
8170 => "100111111100010111101000",
8171 => "100111111100010111101000",
8172 => "011010001000000110011000",
8173 => "000000000000000000000000",
8174 => "000000000000000000000000",
8175 => "010000110100001101000011",
8176 => "010000110100001101000011",
8177 => "000101110001011100010111",
8178 => "000000000000000000000000",
8179 => "001000000010000000100000",
8180 => "011001100110011001100110",
8181 => "011001100110011001100110",
8182 => "010000110100001101000011",
8183 => "010000110100001101000011",
8184 => "000110010001100100011001",
8185 => "000000000000000000000000",
8186 => "000000000000000000000000",
8187 => "000000000000000000000000",
8188 => "000000000000000000000000",
8189 => "000000000000000000000000",
8190 => "000000000000000000000000",
8191 => "000000000000000000000000",
8192 => "000000000000000000000000",
8193 => "000000000000000000000000",
8194 => "000000000000000000000000",
8195 => "000000000000000000000000",
8196 => "000000000000000000000000",
8197 => "000000000000000000000000",
8198 => "000000000000000000000000",
8199 => "000000000000000000000000",
8200 => "000000000000000000000000",
8201 => "000000000000000000000000",
8202 => "000000000000000000000000",
8203 => "000000000000000000000000",
8204 => "000000000000000000000000",
8205 => "000000000000000000000000",
8206 => "000000000000000000000000",
8207 => "000000000000000000000000",
8208 => "000000000000000000000000",
8209 => "000000000000000000000000",
8210 => "000000000000000000000000",
8211 => "000000000000000000000000",
8212 => "000000000000000000000000",
8213 => "000000000000000000000000",
8214 => "000000000000000000000000",
8215 => "000000000000000000000000",
8216 => "000000000000000000000000",
8217 => "000000000000000000000000",
8218 => "000000000000000000000000",
8219 => "000000000000000000000000",
8220 => "000000000000000000000000",
8221 => "000000000000000000000000",
8222 => "000000000000000000000000",
8223 => "000000000000000000000000",
8224 => "000000000000000000000000",
8225 => "000000000000000000000000",
8226 => "000000000000000000000000",
8227 => "000000000000000000000000",
8228 => "000000000000000000000000",
8229 => "000000000000000000000000",
8230 => "000000000000000000000000",
8231 => "000000000000000000000000",
8232 => "000000000000000000000000",
8233 => "000000000000000000000000",
8234 => "000000000000000000000000",
8235 => "000000000000000000000000",
8236 => "000000000000000000000000",
8237 => "000000000000000000000000",
8238 => "000000000000000000000000",
8239 => "000000000000000000000000",
8240 => "000000000000000000000000",
8241 => "000000000000000000000000",
8242 => "000000000000000000000000",
8243 => "000000000000000000000000",
8244 => "000000000000000000000000",
8245 => "000000000000000000000000",
8246 => "000000000000000000000000",
8247 => "000000000000000000000000",
8248 => "000000000000000000000000",
8249 => "000000000000000000000000",
8250 => "000000000000000000000000",
8251 => "000000000000000000000000",
8252 => "000000000000000000000000",
8253 => "000000000000000000000000",
8254 => "000000000000000000000000",
8255 => "000000000000000000000000",
8256 => "000000000000000000000000",
8257 => "000000000000000000000000",
8258 => "000000000000000000000000",
8259 => "000000000000000000000000",
8260 => "000000000000000000000000",
8261 => "000000000000000000000000",
8262 => "000000000000000000000000",
8263 => "000000000000000000000000",
8264 => "000000000000000000000000",
8265 => "000000000000000000000000",
8266 => "000000000000000000000000",
8267 => "000000000000000000000000",
8268 => "000000000000000000000000",
8269 => "000000000000000000000000",
8270 => "000000000000000000000000",
8271 => "000000000000000000000000",
8272 => "000000000000000000000000",
8273 => "000000000000000000000000",
8274 => "000000000000000000000000",
8275 => "000000000000000000000000",
8276 => "000000000000000000000000",
8277 => "000000000000000000000000",
8278 => "000000000000000000000000",
8279 => "000000000000000000000000",
8280 => "000000000000000000000000",
8281 => "000000000000000000000000",
8282 => "000000000000000000000000",
8283 => "000000000000000000000000",
8284 => "000000000000000000000000",
8285 => "000000000000000000000000",
8286 => "000000000000000000000000",
8287 => "000000000000000000000000",
8288 => "000000000000000000000000",
8289 => "000000000000000000000000",
8290 => "000000000000000000000000",
8291 => "000000000000000000000000",
8292 => "000000000000000000000000",
8293 => "000000000000000000000000",
8294 => "000000000000000000000000",
8295 => "000000000000000000000000",
8296 => "000000000000000000000000",
8297 => "000000000000000000000000",
8298 => "000000000000000000000000",
8299 => "000000000000000000000000",
8300 => "000000000000000000000000",
8301 => "000000000000000000000000",
8302 => "000000000000000000000000",
8303 => "000001100000011000000110",
8304 => "010000110100001101000011",
8305 => "010000110100001101000011",
8306 => "010111110101111101011111",
8307 => "011001100110011001100110",
8308 => "001111010011110100111101",
8309 => "000000000000000000000000",
8310 => "000001000000010000000100",
8311 => "010000110100001101000011",
8312 => "010000110100001101000011",
8313 => "000100100001001000010010",
8314 => "000000000000000000000000",
8315 => "001111000100101001010111",
8316 => "100111111100010111101000",
8317 => "100111111100010111101000",
8318 => "100111111100010111101000",
8319 => "100111111100010111101000",
8320 => "100111111100010111101000",
8321 => "100111111100010111101000",
8322 => "011010001000000110011000",
8323 => "000000000000000000000000",
8324 => "000000000000000000000000",
8325 => "010000110100001101000011",
8326 => "010000110100001101000011",
8327 => "000101110001011100010111",
8328 => "000000000000000000000000",
8329 => "001000000010000000100000",
8330 => "011001100110011001100110",
8331 => "011001100110011001100110",
8332 => "010000110100001101000011",
8333 => "010000110100001101000011",
8334 => "000110010001100100011001",
8335 => "000000000000000000000000",
8336 => "000000000000000000000000",
8337 => "000000000000000000000000",
8338 => "000000000000000000000000",
8339 => "000000000000000000000000",
8340 => "000000000000000000000000",
8341 => "000000000000000000000000",
8342 => "000000000000000000000000",
8343 => "000000000000000000000000",
8344 => "000000000000000000000000",
8345 => "000000000000000000000000",
8346 => "000000000000000000000000",
8347 => "000000000000000000000000",
8348 => "000000000000000000000000",
8349 => "000000000000000000000000",
8350 => "000000000000000000000000",
8351 => "000000000000000000000000",
8352 => "000000000000000000000000",
8353 => "000000000000000000000000",
8354 => "000000000000000000000000",
8355 => "000000000000000000000000",
8356 => "000000000000000000000000",
8357 => "000000000000000000000000",
8358 => "000000000000000000000000",
8359 => "000000000000000000000000",
8360 => "000000000000000000000000",
8361 => "000000000000000000000000",
8362 => "000000000000000000000000",
8363 => "000000000000000000000000",
8364 => "000000000000000000000000",
8365 => "000000000000000000000000",
8366 => "000000000000000000000000",
8367 => "000000000000000000000000",
8368 => "000000000000000000000000",
8369 => "000000000000000000000000",
8370 => "000000000000000000000000",
8371 => "000000000000000000000000",
8372 => "000000000000000000000000",
8373 => "000000000000000000000000",
8374 => "000000000000000000000000",
8375 => "000000000000000000000000",
8376 => "000000000000000000000000",
8377 => "000000000000000000000000",
8378 => "000000000000000000000000",
8379 => "000000000000000000000000",
8380 => "000000000000000000000000",
8381 => "000000000000000000000000",
8382 => "000000000000000000000000",
8383 => "000000000000000000000000",
8384 => "000000000000000000000000",
8385 => "000000000000000000000000",
8386 => "000000000000000000000000",
8387 => "000000000000000000000000",
8388 => "000000000000000000000000",
8389 => "000000000000000000000000",
8390 => "000000000000000000000000",
8391 => "000000000000000000000000",
8392 => "000000000000000000000000",
8393 => "000000000000000000000000",
8394 => "000000000000000000000000",
8395 => "000000000000000000000000",
8396 => "000000000000000000000000",
8397 => "000000000000000000000000",
8398 => "000000000000000000000000",
8399 => "000000000000000000000000",
8400 => "000000000000000000000000",
8401 => "000000000000000000000000",
8402 => "000000000000000000000000",
8403 => "000000000000000000000000",
8404 => "000000000000000000000000",
8405 => "000000000000000000000000",
8406 => "000000000000000000000000",
8407 => "000000000000000000000000",
8408 => "000000000000000000000000",
8409 => "000000000000000000000000",
8410 => "000000000000000000000000",
8411 => "000000000000000000000000",
8412 => "000000000000000000000000",
8413 => "000000000000000000000000",
8414 => "000000000000000000000000",
8415 => "000000000000000000000000",
8416 => "000000000000000000000000",
8417 => "000000000000000000000000",
8418 => "000000000000000000000000",
8419 => "000000000000000000000000",
8420 => "000000000000000000000000",
8421 => "000000000000000000000000",
8422 => "000000000000000000000000",
8423 => "000000000000000000000000",
8424 => "000000000000000000000000",
8425 => "000000000000000000000000",
8426 => "000000000000000000000000",
8427 => "000000000000000000000000",
8428 => "000000000000000000000000",
8429 => "000000000000000000000000",
8430 => "000000000000000000000000",
8431 => "000000000000000000000000",
8432 => "000000000000000000000000",
8433 => "000000000000000000000000",
8434 => "000000000000000000000000",
8435 => "000000000000000000000000",
8436 => "000000000000000000000000",
8437 => "000000000000000000000000",
8438 => "000000000000000000000000",
8439 => "000000000000000000000000",
8440 => "000000000000000000000000",
8441 => "000000000000000000000000",
8442 => "000000000000000000000000",
8443 => "000000000000000000000000",
8444 => "000000000000000000000000",
8445 => "000000000000000000000000",
8446 => "000000000000000000000000",
8447 => "000000000000000000000000",
8448 => "000000000000000000000000",
8449 => "000000000000000000000000",
8450 => "000000000000000000000000",
8451 => "000000000000000000000000",
8452 => "000000000000000000000000",
8453 => "000001100000011000000110",
8454 => "010000110100001101000011",
8455 => "010000110100001101000011",
8456 => "010111110101111101011111",
8457 => "011001100110011001100110",
8458 => "001111010011110100111101",
8459 => "000000000000000000000000",
8460 => "000001000000010000000100",
8461 => "010000110100001101000011",
8462 => "010000110100001101000011",
8463 => "000100100001001000010010",
8464 => "000000000000000000000000",
8465 => "001111000100101001010111",
8466 => "100111111100010111101000",
8467 => "100111111100010111101000",
8468 => "100111111100010111101000",
8469 => "100111111100010111101000",
8470 => "100111111100010111101000",
8471 => "100111111100010111101000",
8472 => "011010001000000110011000",
8473 => "000000000000000000000000",
8474 => "000000000000000000000000",
8475 => "010000110100001101000011",
8476 => "010000110100001101000011",
8477 => "000101110001011100010111",
8478 => "000000000000000000000000",
8479 => "001000000010000000100000",
8480 => "011001100110011001100110",
8481 => "011001100110011001100110",
8482 => "010000110100001101000011",
8483 => "010000110100001101000011",
8484 => "000110010001100100011001",
8485 => "000000000000000000000000",
8486 => "000000000000000000000000",
8487 => "000000000000000000000000",
8488 => "000000000000000000000000",
8489 => "000000000000000000000000",
8490 => "000000000000000000000000",
8491 => "000000000000000000000000",
8492 => "000000000000000000000000",
8493 => "000000000000000000000000",
8494 => "000000000000000000000000",
8495 => "000000000000000000000000",
8496 => "000000000000000000000000",
8497 => "000000000000000000000000",
8498 => "000000000000000000000000",
8499 => "000000000000000000000000",
8500 => "000000000000000000000000",
8501 => "000000000000000000000000",
8502 => "000000000000000000000000",
8503 => "000000000000000000000000",
8504 => "000000000000000000000000",
8505 => "000000000000000000000000",
8506 => "000000000000000000000000",
8507 => "000000000000000000000000",
8508 => "000000000000000000000000",
8509 => "000000000000000000000000",
8510 => "000000000000000000000000",
8511 => "000000000000000000000000",
8512 => "000000000000000000000000",
8513 => "000000000000000000000000",
8514 => "000000000000000000000000",
8515 => "000000000000000000000000",
8516 => "000000000000000000000000",
8517 => "000000000000000000000000",
8518 => "000000000000000000000000",
8519 => "000000000000000000000000",
8520 => "000000000000000000000000",
8521 => "000000000000000000000000",
8522 => "000000000000000000000000",
8523 => "000000000000000000000000",
8524 => "000000000000000000000000",
8525 => "000000000000000000000000",
8526 => "000000000000000000000000",
8527 => "000000000000000000000000",
8528 => "000000000000000000000000",
8529 => "000000000000000000000000",
8530 => "000000000000000000000000",
8531 => "000000000000000000000000",
8532 => "000000000000000000000000",
8533 => "000000000000000000000000",
8534 => "000000000000000000000000",
8535 => "000000000000000000000000",
8536 => "000000000000000000000000",
8537 => "000000000000000000000000",
8538 => "000000000000000000000000",
8539 => "000000000000000000000000",
8540 => "000000000000000000000000",
8541 => "000000000000000000000000",
8542 => "000000000000000000000000",
8543 => "000000000000000000000000",
8544 => "000000000000000000000000",
8545 => "000000000000000000000000",
8546 => "000000000000000000000000",
8547 => "000000000000000000000000",
8548 => "000000000000000000000000",
8549 => "000000000000000000000000",
8550 => "000000000000000000000000",
8551 => "000000000000000000000000",
8552 => "000000000000000000000000",
8553 => "000000000000000000000000",
8554 => "000000000000000000000000",
8555 => "000000000000000000000000",
8556 => "000000000000000000000000",
8557 => "000000000000000000000000",
8558 => "000000000000000000000000",
8559 => "000000000000000000000000",
8560 => "000000000000000000000000",
8561 => "000000000000000000000000",
8562 => "000000000000000000000000",
8563 => "000000000000000000000000",
8564 => "000000000000000000000000",
8565 => "000000000000000000000000",
8566 => "000000000000000000000000",
8567 => "000000000000000000000000",
8568 => "000000000000000000000000",
8569 => "000000000000000000000000",
8570 => "000000000000000000000000",
8571 => "000000000000000000000000",
8572 => "000000000000000000000000",
8573 => "000000000000000000000000",
8574 => "000000000000000000000000",
8575 => "000000000000000000000000",
8576 => "000000000000000000000000",
8577 => "000000000000000000000000",
8578 => "000000000000000000000000",
8579 => "000000000000000000000000",
8580 => "000000000000000000000000",
8581 => "000000000000000000000000",
8582 => "000000000000000000000000",
8583 => "000000000000000000000000",
8584 => "000000000000000000000000",
8585 => "000000000000000000000000",
8586 => "000000000000000000000000",
8587 => "000000000000000000000000",
8588 => "000000000000000000000000",
8589 => "000000000000000000000000",
8590 => "000000000000000000000000",
8591 => "000000000000000000000000",
8592 => "000000000000000000000000",
8593 => "000000000000000000000000",
8594 => "000000000000000000000000",
8595 => "000000000000000000000000",
8596 => "000000000000000000000000",
8597 => "000000000000000000000000",
8598 => "000000000000000000000000",
8599 => "000000000000000000000000",
8600 => "000000000000000000000000",
8601 => "000000000000000000000000",
8602 => "000000000000000000000000",
8603 => "000001100000011000000110",
8604 => "010000110100001101000011",
8605 => "010000110100001101000011",
8606 => "010111110101111101011111",
8607 => "011001100110011001100110",
8608 => "001111010011110100111101",
8609 => "000000000000000000000000",
8610 => "000001000000010000000100",
8611 => "010000110100001101000011",
8612 => "010000110100001101000011",
8613 => "000100100001001000010010",
8614 => "000000000000000000000000",
8615 => "001111000100101001010111",
8616 => "100111111100010111101000",
8617 => "100111111100010111101000",
8618 => "100111111100010111101000",
8619 => "100111111100010111101000",
8620 => "100111111100010111101000",
8621 => "100111111100010111101000",
8622 => "011010001000000110011000",
8623 => "000000000000000000000000",
8624 => "000000000000000000000000",
8625 => "010000110100001101000011",
8626 => "010000110100001101000011",
8627 => "000101110001011100010111",
8628 => "000000000000000000000000",
8629 => "001000000010000000100000",
8630 => "011001100110011001100110",
8631 => "011001100110011001100110",
8632 => "010000110100001101000011",
8633 => "010000110100001101000011",
8634 => "000110010001100100011001",
8635 => "000000000000000000000000",
8636 => "000000000000000000000000",
8637 => "000000000000000000000000",
8638 => "000000000000000000000000",
8639 => "000000000000000000000000",
8640 => "000000000000000000000000",
8641 => "000000000000000000000000",
8642 => "000000000000000000000000",
8643 => "000000000000000000000000",
8644 => "000000000000000000000000",
8645 => "000000000000000000000000",
8646 => "000000000000000000000000",
8647 => "000000000000000000000000",
8648 => "000000000000000000000000",
8649 => "000000000000000000000000",
8650 => "000000000000000000000000",
8651 => "000000000000000000000000",
8652 => "000000000000000000000000",
8653 => "000000000000000000000000",
8654 => "000000000000000000000000",
8655 => "000000000000000000000000",
8656 => "000000000000000000000000",
8657 => "000000000000000000000000",
8658 => "000000000000000000000000",
8659 => "000000000000000000000000",
8660 => "000000000000000000000000",
8661 => "000000000000000000000000",
8662 => "000000000000000000000000",
8663 => "000000000000000000000000",
8664 => "000000000000000000000000",
8665 => "000000000000000000000000",
8666 => "000000000000000000000000",
8667 => "000000000000000000000000",
8668 => "000000000000000000000000",
8669 => "000000000000000000000000",
8670 => "000000000000000000000000",
8671 => "000000000000000000000000",
8672 => "000000000000000000000000",
8673 => "000000000000000000000000",
8674 => "000000000000000000000000",
8675 => "000000000000000000000000",
8676 => "000000000000000000000000",
8677 => "000000000000000000000000",
8678 => "000000000000000000000000",
8679 => "000000000000000000000000",
8680 => "000000000000000000000000",
8681 => "000000000000000000000000",
8682 => "000000000000000000000000",
8683 => "000000000000000000000000",
8684 => "000000000000000000000000",
8685 => "000000000000000000000000",
8686 => "000000000000000000000000",
8687 => "000000000000000000000000",
8688 => "000000000000000000000000",
8689 => "000000000000000000000000",
8690 => "000000000000000000000000",
8691 => "000000000000000000000000",
8692 => "000000000000000000000000",
8693 => "000000000000000000000000",
8694 => "000000000000000000000000",
8695 => "000000000000000000000000",
8696 => "000000000000000000000000",
8697 => "000000000000000000000000",
8698 => "000000000000000000000000",
8699 => "000000000000000000000000",
8700 => "000000000000000000000000",
8701 => "000000000000000000000000",
8702 => "000000000000000000000000",
8703 => "000000000000000000000000",
8704 => "000000000000000000000000",
8705 => "000000000000000000000000",
8706 => "000000000000000000000000",
8707 => "000000000000000000000000",
8708 => "000000000000000000000000",
8709 => "000000000000000000000000",
8710 => "000000000000000000000000",
8711 => "000000000000000000000000",
8712 => "000000000000000000000000",
8713 => "000000000000000000000000",
8714 => "000000000000000000000000",
8715 => "000000000000000000000000",
8716 => "000000000000000000000000",
8717 => "000000000000000000000000",
8718 => "000000000000000000000000",
8719 => "000000000000000000000000",
8720 => "000000000000000000000000",
8721 => "000000000000000000000000",
8722 => "000000000000000000000000",
8723 => "000000000000000000000000",
8724 => "000000000000000000000000",
8725 => "000000000000000000000000",
8726 => "000000000000000000000000",
8727 => "000000000000000000000000",
8728 => "000000000000000000000000",
8729 => "000000000000000000000000",
8730 => "000000000000000000000000",
8731 => "000000000000000000000000",
8732 => "000000000000000000000000",
8733 => "000000000000000000000000",
8734 => "000000000000000000000000",
8735 => "000000000000000000000000",
8736 => "000000000000000000000000",
8737 => "000000000000000000000000",
8738 => "000000000000000000000000",
8739 => "000000000000000000000000",
8740 => "000000000000000000000000",
8741 => "000000000000000000000000",
8742 => "000000000000000000000000",
8743 => "000000000000000000000000",
8744 => "000000000000000000000000",
8745 => "000000000000000000000000",
8746 => "000000000000000000000000",
8747 => "000000000000000000000000",
8748 => "000000000000000000000000",
8749 => "000000000000000000000000",
8750 => "000000000000000000000000",
8751 => "000000000000000000000000",
8752 => "000000000000000000000000",
8753 => "000001100000011000000110",
8754 => "010000110100001101000011",
8755 => "010000110100001101000011",
8756 => "010111110101111101011111",
8757 => "011001100110011001100110",
8758 => "001111010011110100111101",
8759 => "000000000000000000000000",
8760 => "000001000000010000000100",
8761 => "010000110100001101000011",
8762 => "010000110100001101000011",
8763 => "000100100001001000010010",
8764 => "000000000000000000000000",
8765 => "001111000100101001010111",
8766 => "100111111100010111101000",
8767 => "100111111100010111101000",
8768 => "100111111100010111101000",
8769 => "100111111100010111101000",
8770 => "100111111100010111101000",
8771 => "100111111100010111101000",
8772 => "011010001000000110011000",
8773 => "000000000000000000000000",
8774 => "000000000000000000000000",
8775 => "010000110100001101000011",
8776 => "010000110100001101000011",
8777 => "000101110001011100010111",
8778 => "000000000000000000000000",
8779 => "001000000010000000100000",
8780 => "011001100110011001100110",
8781 => "011001100110011001100110",
8782 => "010000110100001101000011",
8783 => "010000110100001101000011",
8784 => "000110010001100100011001",
8785 => "000000000000000000000000",
8786 => "000000000000000000000000",
8787 => "000000000000000000000000",
8788 => "000000000000000000000000",
8789 => "000000000000000000000000",
8790 => "000000000000000000000000",
8791 => "000000000000000000000000",
8792 => "000000000000000000000000",
8793 => "000000000000000000000000",
8794 => "000000000000000000000000",
8795 => "000000000000000000000000",
8796 => "000000000000000000000000",
8797 => "000000000000000000000000",
8798 => "000000000000000000000000",
8799 => "000000000000000000000000",
8800 => "000000000000000000000000",
8801 => "000000000000000000000000",
8802 => "000000000000000000000000",
8803 => "000000000000000000000000",
8804 => "000000000000000000000000",
8805 => "000000000000000000000000",
8806 => "000000000000000000000000",
8807 => "000000000000000000000000",
8808 => "000000000000000000000000",
8809 => "000000000000000000000000",
8810 => "000000000000000000000000",
8811 => "000000000000000000000000",
8812 => "000000000000000000000000",
8813 => "000000000000000000000000",
8814 => "000000000000000000000000",
8815 => "000000000000000000000000",
8816 => "000000000000000000000000",
8817 => "000000000000000000000000",
8818 => "000000000000000000000000",
8819 => "000000000000000000000000",
8820 => "000000000000000000000000",
8821 => "000000000000000000000000",
8822 => "000000000000000000000000",
8823 => "000000000000000000000000",
8824 => "000000000000000000000000",
8825 => "000000000000000000000000",
8826 => "000000000000000000000000",
8827 => "000000000000000000000000",
8828 => "000000000000000000000000",
8829 => "000000000000000000000000",
8830 => "000000000000000000000000",
8831 => "000000000000000000000000",
8832 => "000000000000000000000000",
8833 => "000000000000000000000000",
8834 => "000000000000000000000000",
8835 => "000000000000000000000000",
8836 => "000000000000000000000000",
8837 => "000000000000000000000000",
8838 => "000000000000000000000000",
8839 => "000000000000000000000000",
8840 => "000000000000000000000000",
8841 => "000000000000000000000000",
8842 => "000000000000000000000000",
8843 => "000000000000000000000000",
8844 => "000000000000000000000000",
8845 => "000000000000000000000000",
8846 => "000000000000000000000000",
8847 => "000000000000000000000000",
8848 => "000000000000000000000000",
8849 => "000000000000000000000000",
8850 => "000000000000000000000000",
8851 => "000000000000000000000000",
8852 => "000000000000000000000000",
8853 => "000000000000000000000000",
8854 => "000000000000000000000000",
8855 => "000000000000000000000000",
8856 => "000000000000000000000000",
8857 => "000000000000000000000000",
8858 => "000000000000000000000000",
8859 => "000000000000000000000000",
8860 => "000000000000000000000000",
8861 => "000000000000000000000000",
8862 => "000000000000000000000000",
8863 => "000000000000000000000000",
8864 => "000000000000000000000000",
8865 => "000000000000000000000000",
8866 => "000000000000000000000000",
8867 => "000000000000000000000000",
8868 => "000000000000000000000000",
8869 => "000000000000000000000000",
8870 => "000000000000000000000000",
8871 => "000000000000000000000000",
8872 => "000000000000000000000000",
8873 => "000000000000000000000000",
8874 => "000000000000000000000000",
8875 => "000000000000000000000000",
8876 => "000000000000000000000000",
8877 => "000000000000000000000000",
8878 => "000000000000000000000000",
8879 => "000000000000000000000000",
8880 => "000000000000000000000000",
8881 => "000000000000000000000000",
8882 => "000000000000000000000000",
8883 => "000000000000000000000000",
8884 => "000000000000000000000000",
8885 => "000000000000000000000000",
8886 => "000000000000000000000000",
8887 => "000000000000000000000000",
8888 => "000000000000000000000000",
8889 => "000000000000000000000000",
8890 => "000000000000000000000000",
8891 => "000000000000000000000000",
8892 => "000000000000000000000000",
8893 => "000000000000000000000000",
8894 => "000000000000000000000000",
8895 => "000000000000000000000000",
8896 => "000000000000000000000000",
8897 => "000000000000000000000000",
8898 => "000000000000000000000000",
8899 => "000000000000000000000000",
8900 => "000000000000000000000000",
8901 => "000000000000000000000000",
8902 => "000000000000000000000000",
8903 => "000001100000011000000110",
8904 => "010000110100001101000011",
8905 => "010000110100001101000011",
8906 => "010111110101111101011111",
8907 => "011001100110011001100110",
8908 => "001111010011110100111101",
8909 => "000000000000000000000000",
8910 => "000001000000010000000100",
8911 => "010000110100001101000011",
8912 => "010000110100001101000011",
8913 => "000100100001001000010010",
8914 => "000000000000000000000000",
8915 => "001111000100101001010111",
8916 => "100111111100010111101000",
8917 => "100111111100010111101000",
8918 => "100111111100010111101000",
8919 => "100111111100010111101000",
8920 => "100111111100010111101000",
8921 => "100111111100010111101000",
8922 => "011010001000000110011000",
8923 => "000000000000000000000000",
8924 => "000000000000000000000000",
8925 => "010000110100001101000011",
8926 => "010000110100001101000011",
8927 => "000101110001011100010111",
8928 => "000000000000000000000000",
8929 => "001000000010000000100000",
8930 => "011001100110011001100110",
8931 => "011001100110011001100110",
8932 => "010000110100001101000011",
8933 => "010000110100001101000011",
8934 => "000110010001100100011001",
8935 => "000000000000000000000000",
8936 => "000000000000000000000000",
8937 => "000000000000000000000000",
8938 => "000000000000000000000000",
8939 => "000000000000000000000000",
8940 => "000000000000000000000000",
8941 => "000000000000000000000000",
8942 => "000000000000000000000000",
8943 => "000000000000000000000000",
8944 => "000000000000000000000000",
8945 => "000000000000000000000000",
8946 => "000000000000000000000000",
8947 => "000000000000000000000000",
8948 => "000000000000000000000000",
8949 => "000000000000000000000000",
8950 => "000000000000000000000000",
8951 => "000000000000000000000000",
8952 => "000000000000000000000000",
8953 => "000000000000000000000000",
8954 => "000000000000000000000000",
8955 => "000000000000000000000000",
8956 => "000000000000000000000000",
8957 => "000000000000000000000000",
8958 => "000000000000000000000000",
8959 => "000000000000000000000000",
8960 => "000000000000000000000000",
8961 => "000000000000000000000000",
8962 => "000000000000000000000000",
8963 => "000000000000000000000000",
8964 => "000000000000000000000000",
8965 => "000000000000000000000000",
8966 => "000000000000000000000000",
8967 => "000000000000000000000000",
8968 => "000000000000000000000000",
8969 => "000000000000000000000000",
8970 => "000000000000000000000000",
8971 => "000000000000000000000000",
8972 => "000000000000000000000000",
8973 => "000000000000000000000000",
8974 => "000000000000000000000000",
8975 => "000000000000000000000000",
8976 => "000000000000000000000000",
8977 => "000000000000000000000000",
8978 => "000000000000000000000000",
8979 => "000000000000000000000000",
8980 => "000000000000000000000000",
8981 => "000000000000000000000000",
8982 => "000000000000000000000000",
8983 => "000000000000000000000000",
8984 => "000000000000000000000000",
8985 => "000000000000000000000000",
8986 => "000000000000000000000000",
8987 => "000000000000000000000000",
8988 => "000000000000000000000000",
8989 => "000000000000000000000000",
8990 => "000000000000000000000000",
8991 => "000000000000000000000000",
8992 => "000000000000000000000000",
8993 => "000000000000000000000000",
8994 => "000000000000000000000000",
8995 => "000000000000000000000000",
8996 => "000000000000000000000000",
8997 => "000000000000000000000000",
8998 => "000000000000000000000000",
8999 => "000000000000000000000000",
9000 => "000000000000000000000000",
9001 => "000000000000000000000000",
9002 => "000000000000000000000000",
9003 => "000000000000000000000000",
9004 => "000000000000000000000000",
9005 => "000000000000000000000000",
9006 => "000000000000000000000000",
9007 => "000000000000000000000000",
9008 => "000000000000000000000000",
9009 => "000000000000000000000000",
9010 => "000000000000000000000000",
9011 => "000000000000000000000000",
9012 => "000000000000000000000000",
9013 => "000000000000000000000000",
9014 => "000000000000000000000000",
9015 => "000000000000000000000000",
9016 => "000000000000000000000000",
9017 => "000000000000000000000000",
9018 => "000000000000000000000000",
9019 => "000000000000000000000000",
9020 => "000000000000000000000000",
9021 => "000000000000000000000000",
9022 => "000000000000000000000000",
9023 => "000000000000000000000000",
9024 => "000000000000000000000000",
9025 => "000000000000000000000000",
9026 => "000000000000000000000000",
9027 => "000000000000000000000000",
9028 => "000000000000000000000000",
9029 => "000000000000000000000000",
9030 => "000000000000000000000000",
9031 => "000000000000000000000000",
9032 => "000000000000000000000000",
9033 => "000000000000000000000000",
9034 => "000000000000000000000000",
9035 => "000000000000000000000000",
9036 => "000000000000000000000000",
9037 => "000000000000000000000000",
9038 => "000000000000000000000000",
9039 => "000000000000000000000000",
9040 => "000000000000000000000000",
9041 => "000000000000000000000000",
9042 => "000000000000000000000000",
9043 => "000000000000000000000000",
9044 => "000000000000000000000000",
9045 => "000000000000000000000000",
9046 => "000000000000000000000000",
9047 => "000000000000000000000000",
9048 => "000000000000000000000000",
9049 => "000000000000000000000000",
9050 => "000000000000000000000000",
9051 => "000000000000000000000000",
9052 => "000000000000000000000000",
9053 => "000001100000011000000110",
9054 => "010000110100001101000011",
9055 => "010000110100001101000011",
9056 => "010111110101111101011111",
9057 => "011001100110011001100110",
9058 => "001111010011110100111101",
9059 => "000000000000000000000000",
9060 => "000001000000010000000100",
9061 => "010000110100001101000011",
9062 => "010000110100001101000011",
9063 => "000101010001010100010101",
9064 => "000001000000010000000100",
9065 => "001110110100100001010100",
9066 => "100101011011100111011010",
9067 => "100101011011100111011010",
9068 => "100111111100010111101000",
9069 => "100111111100010111101000",
9070 => "100110001011110111011110",
9071 => "100101011011100111011010",
9072 => "011000110111101110010000",
9073 => "000001000000010000000100",
9074 => "000001000000010000000100",
9075 => "010000110100001101000011",
9076 => "010000110100001101000011",
9077 => "000101110001011100010111",
9078 => "000000000000000000000000",
9079 => "001000000010000000100000",
9080 => "011001100110011001100110",
9081 => "011001100110011001100110",
9082 => "010000110100001101000011",
9083 => "010000110100001101000011",
9084 => "000110010001100100011001",
9085 => "000000000000000000000000",
9086 => "000000000000000000000000",
9087 => "000000000000000000000000",
9088 => "000000000000000000000000",
9089 => "000000000000000000000000",
9090 => "000000000000000000000000",
9091 => "000000000000000000000000",
9092 => "000000000000000000000000",
9093 => "000000000000000000000000",
9094 => "000000000000000000000000",
9095 => "000000000000000000000000",
9096 => "000000000000000000000000",
9097 => "000000000000000000000000",
9098 => "000000000000000000000000",
9099 => "000000000000000000000000",
9100 => "000000000000000000000000",
9101 => "000000000000000000000000",
9102 => "000000000000000000000000",
9103 => "000000000000000000000000",
9104 => "000000000000000000000000",
9105 => "000000000000000000000000",
9106 => "000000000000000000000000",
9107 => "000000000000000000000000",
9108 => "000000000000000000000000",
9109 => "000000000000000000000000",
9110 => "000000000000000000000000",
9111 => "000000000000000000000000",
9112 => "000000000000000000000000",
9113 => "000000000000000000000000",
9114 => "000000000000000000000000",
9115 => "000000000000000000000000",
9116 => "000000000000000000000000",
9117 => "000000000000000000000000",
9118 => "000000000000000000000000",
9119 => "000000000000000000000000",
9120 => "000000000000000000000000",
9121 => "000000000000000000000000",
9122 => "000000000000000000000000",
9123 => "000000000000000000000000",
9124 => "000000000000000000000000",
9125 => "000000000000000000000000",
9126 => "000000000000000000000000",
9127 => "000000000000000000000000",
9128 => "000000000000000000000000",
9129 => "000000000000000000000000",
9130 => "000000000000000000000000",
9131 => "000000000000000000000000",
9132 => "000000000000000000000000",
9133 => "000000000000000000000000",
9134 => "000000000000000000000000",
9135 => "000000000000000000000000",
9136 => "000000000000000000000000",
9137 => "000000000000000000000000",
9138 => "000000000000000000000000",
9139 => "000000000000000000000000",
9140 => "000000000000000000000000",
9141 => "000000000000000000000000",
9142 => "000000000000000000000000",
9143 => "000000000000000000000000",
9144 => "000000000000000000000000",
9145 => "000000000000000000000000",
9146 => "000000000000000000000000",
9147 => "000000000000000000000000",
9148 => "000000000000000000000000",
9149 => "000000000000000000000000",
9150 => "000000000000000000000000",
9151 => "000000000000000000000000",
9152 => "000000000000000000000000",
9153 => "000000000000000000000000",
9154 => "000000000000000000000000",
9155 => "000000000000000000000000",
9156 => "000000000000000000000000",
9157 => "000000000000000000000000",
9158 => "000000000000000000000000",
9159 => "000000000000000000000000",
9160 => "000000000000000000000000",
9161 => "000000000000000000000000",
9162 => "000000000000000000000000",
9163 => "000000000000000000000000",
9164 => "000000000000000000000000",
9165 => "000000000000000000000000",
9166 => "000000000000000000000000",
9167 => "000000000000000000000000",
9168 => "000000000000000000000000",
9169 => "000000000000000000000000",
9170 => "000000000000000000000000",
9171 => "000000000000000000000000",
9172 => "000000000000000000000000",
9173 => "000000000000000000000000",
9174 => "000000000000000000000000",
9175 => "000000000000000000000000",
9176 => "000000000000000000000000",
9177 => "000000000000000000000000",
9178 => "000000000000000000000000",
9179 => "000000000000000000000000",
9180 => "000000000000000000000000",
9181 => "000000000000000000000000",
9182 => "000000000000000000000000",
9183 => "000000000000000000000000",
9184 => "000000000000000000000000",
9185 => "000000000000000000000000",
9186 => "000000000000000000000000",
9187 => "000000000000000000000000",
9188 => "000000000000000000000000",
9189 => "000000000000000000000000",
9190 => "000000000000000000000000",
9191 => "000000000000000000000000",
9192 => "000000000000000000000000",
9193 => "000000000000000000000000",
9194 => "000000000000000000000000",
9195 => "000000000000000000000000",
9196 => "000000000000000000000000",
9197 => "000000000000000000000000",
9198 => "000000000000000000000000",
9199 => "000000000000000000000000",
9200 => "000000000000000000000000",
9201 => "000000000000000000000000",
9202 => "000000000000000000000000",
9203 => "000001100000011000000110",
9204 => "010000110100001101000011",
9205 => "010000110100001101000011",
9206 => "010111110101111101011111",
9207 => "011001100110011001100110",
9208 => "001111010011110100111101",
9209 => "000000000000000000000000",
9210 => "000001000000010000000100",
9211 => "010000110100001101000011",
9212 => "010000110100001101000011",
9213 => "010000110100001101000011",
9214 => "010000110100001101000011",
9215 => "001010100010101000101010",
9216 => "000000000000000000000000",
9217 => "000001010000011000000111",
9218 => "100111111100010111101000",
9219 => "100111111100010111101000",
9220 => "001100100011111001001001",
9221 => "000000000000000000000000",
9222 => "000101110001011100010111",
9223 => "010000110100001101000011",
9224 => "010000110100001101000011",
9225 => "010000110100001101000011",
9226 => "010000110100001101000011",
9227 => "000101110001011100010111",
9228 => "000000000000000000000000",
9229 => "001000000010000000100000",
9230 => "011001100110011001100110",
9231 => "011001100110011001100110",
9232 => "010000110100001101000011",
9233 => "010000110100001101000011",
9234 => "000110010001100100011001",
9235 => "000000000000000000000000",
9236 => "000000000000000000000000",
9237 => "000000000000000000000000",
9238 => "000000000000000000000000",
9239 => "000000000000000000000000",
9240 => "000000000000000000000000",
9241 => "000000000000000000000000",
9242 => "000000000000000000000000",
9243 => "000000000000000000000000",
9244 => "000000000000000000000000",
9245 => "000000000000000000000000",
9246 => "000000000000000000000000",
9247 => "000000000000000000000000",
9248 => "000000000000000000000000",
9249 => "000000000000000000000000",
9250 => "000000000000000000000000",
9251 => "000000000000000000000000",
9252 => "000000000000000000000000",
9253 => "000000000000000000000000",
9254 => "000000000000000000000000",
9255 => "000000000000000000000000",
9256 => "000000000000000000000000",
9257 => "000000000000000000000000",
9258 => "000000000000000000000000",
9259 => "000000000000000000000000",
9260 => "000000000000000000000000",
9261 => "000000000000000000000000",
9262 => "000000000000000000000000",
9263 => "000000000000000000000000",
9264 => "000000000000000000000000",
9265 => "000000000000000000000000",
9266 => "000000000000000000000000",
9267 => "000000000000000000000000",
9268 => "000000000000000000000000",
9269 => "000000000000000000000000",
9270 => "000000000000000000000000",
9271 => "000000000000000000000000",
9272 => "000000000000000000000000",
9273 => "000000000000000000000000",
9274 => "000000000000000000000000",
9275 => "000000000000000000000000",
9276 => "000000000000000000000000",
9277 => "000000000000000000000000",
9278 => "000000000000000000000000",
9279 => "000000000000000000000000",
9280 => "000000000000000000000000",
9281 => "000000000000000000000000",
9282 => "000000000000000000000000",
9283 => "000000000000000000000000",
9284 => "000000000000000000000000",
9285 => "000000000000000000000000",
9286 => "000000000000000000000000",
9287 => "000000000000000000000000",
9288 => "000000000000000000000000",
9289 => "000000000000000000000000",
9290 => "000000000000000000000000",
9291 => "000000000000000000000000",
9292 => "000000000000000000000000",
9293 => "000000000000000000000000",
9294 => "000000000000000000000000",
9295 => "000000000000000000000000",
9296 => "000000000000000000000000",
9297 => "000000000000000000000000",
9298 => "000000000000000000000000",
9299 => "000000000000000000000000",
9300 => "000000000000000000000000",
9301 => "000000000000000000000000",
9302 => "000000000000000000000000",
9303 => "000000000000000000000000",
9304 => "000000000000000000000000",
9305 => "000000000000000000000000",
9306 => "000000000000000000000000",
9307 => "000000000000000000000000",
9308 => "000000000000000000000000",
9309 => "000000000000000000000000",
9310 => "000000000000000000000000",
9311 => "000000000000000000000000",
9312 => "000000000000000000000000",
9313 => "000000000000000000000000",
9314 => "000000000000000000000000",
9315 => "000000000000000000000000",
9316 => "000000000000000000000000",
9317 => "000000000000000000000000",
9318 => "000000000000000000000000",
9319 => "000000000000000000000000",
9320 => "000000000000000000000000",
9321 => "000000000000000000000000",
9322 => "000000000000000000000000",
9323 => "000000000000000000000000",
9324 => "000000000000000000000000",
9325 => "000000000000000000000000",
9326 => "000000000000000000000000",
9327 => "000000000000000000000000",
9328 => "000000000000000000000000",
9329 => "000000000000000000000000",
9330 => "000000000000000000000000",
9331 => "000000000000000000000000",
9332 => "000000000000000000000000",
9333 => "000000000000000000000000",
9334 => "000000000000000000000000",
9335 => "000000000000000000000000",
9336 => "000000000000000000000000",
9337 => "000000000000000000000000",
9338 => "000000000000000000000000",
9339 => "000000000000000000000000",
9340 => "000000000000000000000000",
9341 => "000000000000000000000000",
9342 => "000000000000000000000000",
9343 => "000000000000000000000000",
9344 => "000000000000000000000000",
9345 => "000000000000000000000000",
9346 => "000000000000000000000000",
9347 => "000000000000000000000000",
9348 => "000000000000000000000000",
9349 => "000000000000000000000000",
9350 => "000000000000000000000000",
9351 => "000000000000000000000000",
9352 => "000000000000000000000000",
9353 => "000001100000011000000110",
9354 => "010000110100001101000011",
9355 => "010000110100001101000011",
9356 => "010111110101111101011111",
9357 => "011001100110011001100110",
9358 => "001111010011110100111101",
9359 => "000000000000000000000000",
9360 => "000001000000010000000100",
9361 => "010000110100001101000011",
9362 => "010000110100001101000011",
9363 => "010000110100001101000011",
9364 => "010000110100001101000011",
9365 => "001010100010101000101010",
9366 => "000000000000000000000000",
9367 => "000001010000011000000111",
9368 => "100111111100010111101000",
9369 => "100111111100010111101000",
9370 => "001100100011111001001001",
9371 => "000000000000000000000000",
9372 => "000101110001011100010111",
9373 => "010000110100001101000011",
9374 => "010000110100001101000011",
9375 => "010000110100001101000011",
9376 => "010000110100001101000011",
9377 => "000101110001011100010111",
9378 => "000000000000000000000000",
9379 => "001000000010000000100000",
9380 => "011001100110011001100110",
9381 => "011001100110011001100110",
9382 => "010000110100001101000011",
9383 => "010000110100001101000011",
9384 => "000110010001100100011001",
9385 => "000000000000000000000000",
9386 => "000000000000000000000000",
9387 => "000000000000000000000000",
9388 => "000000000000000000000000",
9389 => "000000000000000000000000",
9390 => "000000000000000000000000",
9391 => "000000000000000000000000",
9392 => "000000000000000000000000",
9393 => "000000000000000000000000",
9394 => "000000000000000000000000",
9395 => "000000000000000000000000",
9396 => "000000000000000000000000",
9397 => "000000000000000000000000",
9398 => "000000000000000000000000",
9399 => "000000000000000000000000",
9400 => "000000000000000000000000",
9401 => "000000000000000000000000",
9402 => "000000000000000000000000",
9403 => "000000000000000000000000",
9404 => "000000000000000000000000",
9405 => "000000000000000000000000",
9406 => "000000000000000000000000",
9407 => "000000000000000000000000",
9408 => "000000000000000000000000",
9409 => "000000000000000000000000",
9410 => "000000000000000000000000",
9411 => "000000000000000000000000",
9412 => "000000000000000000000000",
9413 => "000000000000000000000000",
9414 => "000000000000000000000000",
9415 => "000000000000000000000000",
9416 => "000000000000000000000000",
9417 => "000000000000000000000000",
9418 => "000000000000000000000000",
9419 => "000000000000000000000000",
9420 => "000000000000000000000000",
9421 => "000000000000000000000000",
9422 => "000000000000000000000000",
9423 => "000000000000000000000000",
9424 => "000000000000000000000000",
9425 => "000000000000000000000000",
9426 => "000000000000000000000000",
9427 => "000000000000000000000000",
9428 => "000000000000000000000000",
9429 => "000000000000000000000000",
9430 => "000000000000000000000000",
9431 => "000000000000000000000000",
9432 => "000000000000000000000000",
9433 => "000000000000000000000000",
9434 => "000000000000000000000000",
9435 => "000000000000000000000000",
9436 => "000000000000000000000000",
9437 => "000000000000000000000000",
9438 => "000000000000000000000000",
9439 => "000000000000000000000000",
9440 => "000000000000000000000000",
9441 => "000000000000000000000000",
9442 => "000000000000000000000000",
9443 => "000000000000000000000000",
9444 => "000000000000000000000000",
9445 => "000000000000000000000000",
9446 => "000000000000000000000000",
9447 => "000000000000000000000000",
9448 => "000000000000000000000000",
9449 => "000000000000000000000000",
9450 => "000000000000000000000000",
9451 => "000000000000000000000000",
9452 => "000000000000000000000000",
9453 => "000000000000000000000000",
9454 => "000000000000000000000000",
9455 => "000000000000000000000000",
9456 => "000000000000000000000000",
9457 => "000000000000000000000000",
9458 => "000000000000000000000000",
9459 => "000000000000000000000000",
9460 => "000000000000000000000000",
9461 => "000000000000000000000000",
9462 => "000000000000000000000000",
9463 => "000000000000000000000000",
9464 => "000000000000000000000000",
9465 => "000000000000000000000000",
9466 => "000000000000000000000000",
9467 => "000000000000000000000000",
9468 => "000000000000000000000000",
9469 => "000000000000000000000000",
9470 => "000000000000000000000000",
9471 => "000000000000000000000000",
9472 => "000000000000000000000000",
9473 => "000000000000000000000000",
9474 => "000000000000000000000000",
9475 => "000000000000000000000000",
9476 => "000000000000000000000000",
9477 => "000000000000000000000000",
9478 => "000000000000000000000000",
9479 => "000000000000000000000000",
9480 => "000000000000000000000000",
9481 => "000000000000000000000000",
9482 => "000000000000000000000000",
9483 => "000000000000000000000000",
9484 => "000000000000000000000000",
9485 => "000000000000000000000000",
9486 => "000000000000000000000000",
9487 => "000000000000000000000000",
9488 => "000000000000000000000000",
9489 => "000000000000000000000000",
9490 => "000000000000000000000000",
9491 => "000000000000000000000000",
9492 => "000000000000000000000000",
9493 => "000000000000000000000000",
9494 => "000000000000000000000000",
9495 => "000000000000000000000000",
9496 => "000000000000000000000000",
9497 => "000000000000000000000000",
9498 => "000000000000000000000000",
9499 => "000000000000000000000000",
9500 => "000000000000000000000000",
9501 => "000000000000000000000000",
9502 => "000000000000000000000000",
9503 => "000001100000011000000110",
9504 => "010000110100001101000011",
9505 => "010000110100001101000011",
9506 => "010111110101111101011111",
9507 => "011001100110011001100110",
9508 => "001111010011110100111101",
9509 => "000000000000000000000000",
9510 => "000001000000010000000100",
9511 => "010000110100001101000011",
9512 => "010000110100001101000011",
9513 => "010000110100001101000011",
9514 => "010000110100001101000011",
9515 => "001010100010101000101010",
9516 => "000000000000000000000000",
9517 => "000000010000001000000010",
9518 => "001010110011010100111111",
9519 => "001010110011010100111111",
9520 => "000011010001000100010100",
9521 => "000000000000000000000000",
9522 => "000101110001011100010111",
9523 => "010000110100001101000011",
9524 => "010000110100001101000011",
9525 => "010000110100001101000011",
9526 => "010000110100001101000011",
9527 => "000101110001011100010111",
9528 => "000000000000000000000000",
9529 => "001000000010000000100000",
9530 => "011001100110011001100110",
9531 => "011001100110011001100110",
9532 => "010000110100001101000011",
9533 => "010000110100001101000011",
9534 => "000110010001100100011001",
9535 => "000000000000000000000000",
9536 => "000000000000000000000000",
9537 => "000000000000000000000000",
9538 => "000000000000000000000000",
9539 => "000000000000000000000000",
9540 => "000000000000000000000000",
9541 => "000000000000000000000000",
9542 => "000000000000000000000000",
9543 => "000000000000000000000000",
9544 => "000000000000000000000000",
9545 => "000000000000000000000000",
9546 => "000000000000000000000000",
9547 => "000000000000000000000000",
9548 => "000000000000000000000000",
9549 => "000000000000000000000000",
9550 => "000000000000000000000000",
9551 => "000000000000000000000000",
9552 => "000000000000000000000000",
9553 => "000000000000000000000000",
9554 => "000000000000000000000000",
9555 => "000000000000000000000000",
9556 => "000000000000000000000000",
9557 => "000000000000000000000000",
9558 => "000000000000000000000000",
9559 => "000000000000000000000000",
9560 => "000000000000000000000000",
9561 => "000000000000000000000000",
9562 => "000000000000000000000000",
9563 => "000000000000000000000000",
9564 => "000000000000000000000000",
9565 => "000000000000000000000000",
9566 => "000000000000000000000000",
9567 => "000000000000000000000000",
9568 => "000000000000000000000000",
9569 => "000000000000000000000000",
9570 => "000000000000000000000000",
9571 => "000000000000000000000000",
9572 => "000000000000000000000000",
9573 => "000000000000000000000000",
9574 => "000000000000000000000000",
9575 => "000000000000000000000000",
9576 => "000000000000000000000000",
9577 => "000000000000000000000000",
9578 => "000000000000000000000000",
9579 => "000000000000000000000000",
9580 => "000000000000000000000000",
9581 => "000000000000000000000000",
9582 => "000000000000000000000000",
9583 => "000000000000000000000000",
9584 => "000000000000000000000000",
9585 => "000000000000000000000000",
9586 => "000000000000000000000000",
9587 => "000000000000000000000000",
9588 => "000000000000000000000000",
9589 => "000000000000000000000000",
9590 => "000000000000000000000000",
9591 => "000000000000000000000000",
9592 => "000000000000000000000000",
9593 => "000000000000000000000000",
9594 => "000000000000000000000000",
9595 => "000000000000000000000000",
9596 => "000000000000000000000000",
9597 => "000000000000000000000000",
9598 => "000000000000000000000000",
9599 => "000000000000000000000000",
9600 => "000000000000000000000000",
9601 => "000000000000000000000000",
9602 => "000000000000000000000000",
9603 => "000000000000000000000000",
9604 => "000000000000000000000000",
9605 => "000000000000000000000000",
9606 => "000000000000000000000000",
9607 => "000000000000000000000000",
9608 => "000000000000000000000000",
9609 => "000000000000000000000000",
9610 => "000000000000000000000000",
9611 => "000000000000000000000000",
9612 => "000000000000000000000000",
9613 => "000000000000000000000000",
9614 => "000000000000000000000000",
9615 => "000000000000000000000000",
9616 => "000000000000000000000000",
9617 => "000000000000000000000000",
9618 => "000000000000000000000000",
9619 => "000000000000000000000000",
9620 => "000000000000000000000000",
9621 => "000000000000000000000000",
9622 => "000000000000000000000000",
9623 => "000000000000000000000000",
9624 => "000000000000000000000000",
9625 => "000000000000000000000000",
9626 => "000000000000000000000000",
9627 => "000000000000000000000000",
9628 => "000000000000000000000000",
9629 => "000000000000000000000000",
9630 => "000000000000000000000000",
9631 => "000000000000000000000000",
9632 => "000000000000000000000000",
9633 => "000000000000000000000000",
9634 => "000000000000000000000000",
9635 => "000000000000000000000000",
9636 => "000000000000000000000000",
9637 => "000000000000000000000000",
9638 => "000000000000000000000000",
9639 => "000000000000000000000000",
9640 => "000000000000000000000000",
9641 => "000000000000000000000000",
9642 => "000000000000000000000000",
9643 => "000000000000000000000000",
9644 => "000000000000000000000000",
9645 => "000000000000000000000000",
9646 => "000000000000000000000000",
9647 => "000000000000000000000000",
9648 => "000000000000000000000000",
9649 => "000000000000000000000000",
9650 => "000000000000000000000000",
9651 => "000000000000000000000000",
9652 => "000000000000000000000000",
9653 => "000001100000011000000110",
9654 => "010000110100001101000011",
9655 => "010000110100001101000011",
9656 => "010111110101111101011111",
9657 => "011001100110011001100110",
9658 => "001111010011110100111101",
9659 => "000000000000000000000000",
9660 => "000001000000010000000100",
9661 => "010000110100001101000011",
9662 => "010000110100001101000011",
9663 => "010000110100001101000011",
9664 => "010000110100001101000011",
9665 => "001010100010101000101010",
9666 => "000000000000000000000000",
9667 => "000000000000000000000000",
9668 => "000000000000000000000000",
9669 => "000000000000000000000000",
9670 => "000000000000000000000000",
9671 => "000000000000000000000000",
9672 => "000101110001011100010111",
9673 => "010000110100001101000011",
9674 => "010000110100001101000011",
9675 => "010000110100001101000011",
9676 => "010000110100001101000011",
9677 => "000101110001011100010111",
9678 => "000000000000000000000000",
9679 => "001000000010000000100000",
9680 => "011001100110011001100110",
9681 => "011001100110011001100110",
9682 => "010000110100001101000011",
9683 => "010000110100001101000011",
9684 => "000110010001100100011001",
9685 => "000000000000000000000000",
9686 => "000000000000000000000000",
9687 => "000000000000000000000000",
9688 => "000000000000000000000000",
9689 => "000000000000000000000000",
9690 => "000000000000000000000000",
9691 => "000000000000000000000000",
9692 => "000000000000000000000000",
9693 => "000000000000000000000000",
9694 => "000000000000000000000000",
9695 => "000000000000000000000000",
9696 => "000000000000000000000000",
9697 => "000000000000000000000000",
9698 => "000000000000000000000000",
9699 => "000000000000000000000000",
9700 => "000000000000000000000000",
9701 => "000000000000000000000000",
9702 => "000000000000000000000000",
9703 => "000000000000000000000000",
9704 => "000000000000000000000000",
9705 => "000000000000000000000000",
9706 => "000000000000000000000000",
9707 => "000000000000000000000000",
9708 => "000000000000000000000000",
9709 => "000000000000000000000000",
9710 => "000000000000000000000000",
9711 => "000000000000000000000000",
9712 => "000000000000000000000000",
9713 => "000000000000000000000000",
9714 => "000000000000000000000000",
9715 => "000000000000000000000000",
9716 => "000000000000000000000000",
9717 => "000000000000000000000000",
9718 => "000000000000000000000000",
9719 => "000000000000000000000000",
9720 => "000000000000000000000000",
9721 => "000000000000000000000000",
9722 => "000000000000000000000000",
9723 => "000000000000000000000000",
9724 => "000000000000000000000000",
9725 => "000000000000000000000000",
9726 => "000000000000000000000000",
9727 => "000000000000000000000000",
9728 => "000000000000000000000000",
9729 => "000000000000000000000000",
9730 => "000000000000000000000000",
9731 => "000000000000000000000000",
9732 => "000000000000000000000000",
9733 => "000000000000000000000000",
9734 => "000000000000000000000000",
9735 => "000000000000000000000000",
9736 => "000000000000000000000000",
9737 => "000000000000000000000000",
9738 => "000000000000000000000000",
9739 => "000000000000000000000000",
9740 => "000000000000000000000000",
9741 => "000000000000000000000000",
9742 => "000000000000000000000000",
9743 => "000000000000000000000000",
9744 => "000000000000000000000000",
9745 => "000000000000000000000000",
9746 => "000000000000000000000000",
9747 => "000000000000000000000000",
9748 => "000000000000000000000000",
9749 => "000000000000000000000000",
9750 => "000000000000000000000000",
9751 => "000000000000000000000000",
9752 => "000000000000000000000000",
9753 => "000000000000000000000000",
9754 => "000000000000000000000000",
9755 => "000000000000000000000000",
9756 => "000000000000000000000000",
9757 => "000000000000000000000000",
9758 => "000000000000000000000000",
9759 => "000000000000000000000000",
9760 => "000000000000000000000000",
9761 => "000000000000000000000000",
9762 => "000000000000000000000000",
9763 => "000000000000000000000000",
9764 => "000000000000000000000000",
9765 => "000000000000000000000000",
9766 => "000000000000000000000000",
9767 => "000000000000000000000000",
9768 => "000000000000000000000000",
9769 => "000000000000000000000000",
9770 => "000000000000000000000000",
9771 => "000000000000000000000000",
9772 => "000000000000000000000000",
9773 => "000000000000000000000000",
9774 => "000000000000000000000000",
9775 => "000000000000000000000000",
9776 => "000000000000000000000000",
9777 => "000000000000000000000000",
9778 => "000000000000000000000000",
9779 => "000000000000000000000000",
9780 => "000000000000000000000000",
9781 => "000000000000000000000000",
9782 => "000000000000000000000000",
9783 => "000000000000000000000000",
9784 => "000000000000000000000000",
9785 => "000000000000000000000000",
9786 => "000000000000000000000000",
9787 => "000000000000000000000000",
9788 => "000000000000000000000000",
9789 => "000000000000000000000000",
9790 => "000000000000000000000000",
9791 => "000000000000000000000000",
9792 => "000000000000000000000000",
9793 => "000000000000000000000000",
9794 => "000000000000000000000000",
9795 => "000000000000000000000000",
9796 => "000000000000000000000000",
9797 => "000000000000000000000000",
9798 => "000000000000000000000000",
9799 => "000000000000000000000000",
9800 => "000000000000000000000000",
9801 => "000000000000000000000000",
9802 => "000000000000000000000000",
9803 => "000001100000011000000110",
9804 => "010000110100001101000011",
9805 => "010000110100001101000011",
9806 => "010111110101111101011111",
9807 => "011001100110011001100110",
9808 => "001111010011110100111101",
9809 => "000000000000000000000000",
9810 => "000001000000010000000100",
9811 => "010000110100001101000011",
9812 => "010000110100001101000011",
9813 => "010000110100001101000011",
9814 => "010000110100001101000011",
9815 => "001100110011001100110011",
9816 => "000110010001100100011001",
9817 => "000110010001100100011001",
9818 => "000110010001100100011001",
9819 => "000110010001100100011001",
9820 => "000110010001100100011001",
9821 => "000110010001100100011001",
9822 => "001010000010100000101000",
9823 => "010000110100001101000011",
9824 => "010000110100001101000011",
9825 => "010000110100001101000011",
9826 => "010000110100001101000011",
9827 => "000101110001011100010111",
9828 => "000000000000000000000000",
9829 => "001000000010000000100000",
9830 => "011001100110011001100110",
9831 => "011001100110011001100110",
9832 => "010000110100001101000011",
9833 => "010000110100001101000011",
9834 => "000110010001100100011001",
9835 => "000000000000000000000000",
9836 => "000000000000000000000000",
9837 => "000000000000000000000000",
9838 => "000000000000000000000000",
9839 => "000000000000000000000000",
9840 => "000000000000000000000000",
9841 => "000000000000000000000000",
9842 => "000000000000000000000000",
9843 => "000000000000000000000000",
9844 => "000000000000000000000000",
9845 => "000000000000000000000000",
9846 => "000000000000000000000000",
9847 => "000000000000000000000000",
9848 => "000000000000000000000000",
9849 => "000000000000000000000000",
9850 => "000000000000000000000000",
9851 => "000000000000000000000000",
9852 => "000000000000000000000000",
9853 => "000000000000000000000000",
9854 => "000000000000000000000000",
9855 => "000000000000000000000000",
9856 => "000000000000000000000000",
9857 => "000000000000000000000000",
9858 => "000000000000000000000000",
9859 => "000000000000000000000000",
9860 => "000000000000000000000000",
9861 => "000000000000000000000000",
9862 => "000000000000000000000000",
9863 => "000000000000000000000000",
9864 => "000000000000000000000000",
9865 => "000000000000000000000000",
9866 => "000000000000000000000000",
9867 => "000000000000000000000000",
9868 => "000000000000000000000000",
9869 => "000000000000000000000000",
9870 => "000000000000000000000000",
9871 => "000000000000000000000000",
9872 => "000000000000000000000000",
9873 => "000000000000000000000000",
9874 => "000000000000000000000000",
9875 => "000000000000000000000000",
9876 => "000000000000000000000000",
9877 => "000000000000000000000000",
9878 => "000000000000000000000000",
9879 => "000000000000000000000000",
9880 => "000000000000000000000000",
9881 => "000000000000000000000000",
9882 => "000000000000000000000000",
9883 => "000000000000000000000000",
9884 => "000000000000000000000000",
9885 => "000000000000000000000000",
9886 => "000000000000000000000000",
9887 => "000000000000000000000000",
9888 => "000000000000000000000000",
9889 => "000000000000000000000000",
9890 => "000000000000000000000000",
9891 => "000000000000000000000000",
9892 => "000000000000000000000000",
9893 => "000000000000000000000000",
9894 => "000000000000000000000000",
9895 => "000000000000000000000000",
9896 => "000000000000000000000000",
9897 => "000000000000000000000000",
9898 => "000000000000000000000000",
9899 => "000000000000000000000000",
9900 => "000000000000000000000000",
9901 => "000000000000000000000000",
9902 => "000000000000000000000000",
9903 => "000000000000000000000000",
9904 => "000000000000000000000000",
9905 => "000000000000000000000000",
9906 => "000000000000000000000000",
9907 => "000000000000000000000000",
9908 => "000000000000000000000000",
9909 => "000000000000000000000000",
9910 => "000000000000000000000000",
9911 => "000000000000000000000000",
9912 => "000000000000000000000000",
9913 => "000000000000000000000000",
9914 => "000000000000000000000000",
9915 => "000000000000000000000000",
9916 => "000000000000000000000000",
9917 => "000000000000000000000000",
9918 => "000000000000000000000000",
9919 => "000000000000000000000000",
9920 => "000000000000000000000000",
9921 => "000000000000000000000000",
9922 => "000000000000000000000000",
9923 => "000000000000000000000000",
9924 => "000000000000000000000000",
9925 => "000000000000000000000000",
9926 => "000000000000000000000000",
9927 => "000000000000000000000000",
9928 => "000000000000000000000000",
9929 => "000000000000000000000000",
9930 => "000000000000000000000000",
9931 => "000000000000000000000000",
9932 => "000000000000000000000000",
9933 => "000000000000000000000000",
9934 => "000000000000000000000000",
9935 => "000000000000000000000000",
9936 => "000000000000000000000000",
9937 => "000000000000000000000000",
9938 => "000000000000000000000000",
9939 => "000000000000000000000000",
9940 => "000000000000000000000000",
9941 => "000000000000000000000000",
9942 => "000000000000000000000000",
9943 => "000000000000000000000000",
9944 => "000000000000000000000000",
9945 => "000000000000000000000000",
9946 => "000000000000000000000000",
9947 => "000000000000000000000000",
9948 => "000000000000000000000000",
9949 => "000000000000000000000000",
9950 => "000000000000000000000000",
9951 => "000000000000000000000000",
9952 => "000000000000000000000000",
9953 => "000001100000011000000110",
9954 => "010000110100001101000011",
9955 => "010000110100001101000011",
9956 => "010111110101111101011111",
9957 => "011001100110011001100110",
9958 => "001111010011110100111101",
9959 => "000000000000000000000000",
9960 => "000001000000010000000100",
9961 => "010000110100001101000011",
9962 => "010000110100001101000011",
9963 => "010000110100001101000011",
9964 => "010000110100001101000011",
9965 => "010000110100001101000011",
9966 => "010000110100001101000011",
9967 => "010000110100001101000011",
9968 => "010000110100001101000011",
9969 => "010000110100001101000011",
9970 => "010000110100001101000011",
9971 => "010000110100001101000011",
9972 => "010000110100001101000011",
9973 => "010000110100001101000011",
9974 => "010000110100001101000011",
9975 => "010000110100001101000011",
9976 => "010000110100001101000011",
9977 => "000101110001011100010111",
9978 => "000000000000000000000000",
9979 => "001000000010000000100000",
9980 => "011001100110011001100110",
9981 => "011001100110011001100110",
9982 => "010000110100001101000011",
9983 => "010000110100001101000011",
9984 => "000110010001100100011001",
9985 => "000000000000000000000000",
9986 => "000000000000000000000000",
9987 => "000000000000000000000000",
9988 => "000000000000000000000000",
9989 => "000000000000000000000000",
9990 => "000000000000000000000000",
9991 => "000000000000000000000000",
9992 => "000000000000000000000000",
9993 => "000000000000000000000000",
9994 => "000000000000000000000000",
9995 => "000000000000000000000000",
9996 => "000000000000000000000000",
9997 => "000000000000000000000000",
9998 => "000000000000000000000000",
9999 => "000000000000000000000000",
10000 => "000000000000000000000000",
10001 => "000000000000000000000000",
10002 => "000000000000000000000000",
10003 => "000000000000000000000000",
10004 => "000000000000000000000000",
10005 => "000000000000000000000000",
10006 => "000000000000000000000000",
10007 => "000000000000000000000000",
10008 => "000000000000000000000000",
10009 => "000000000000000000000000",
10010 => "000000000000000000000000",
10011 => "000000000000000000000000",
10012 => "000000000000000000000000",
10013 => "000000000000000000000000",
10014 => "000000000000000000000000",
10015 => "000000000000000000000000",
10016 => "000000000000000000000000",
10017 => "000000000000000000000000",
10018 => "000000000000000000000000",
10019 => "000000000000000000000000",
10020 => "000000000000000000000000",
10021 => "000000000000000000000000",
10022 => "000000000000000000000000",
10023 => "000000000000000000000000",
10024 => "000000000000000000000000",
10025 => "000000000000000000000000",
10026 => "000000000000000000000000",
10027 => "000000000000000000000000",
10028 => "000000000000000000000000",
10029 => "000000000000000000000000",
10030 => "000000000000000000000000",
10031 => "000000000000000000000000",
10032 => "000000000000000000000000",
10033 => "000000000000000000000000",
10034 => "000000000000000000000000",
10035 => "000000000000000000000000",
10036 => "000000000000000000000000",
10037 => "000000000000000000000000",
10038 => "000000000000000000000000",
10039 => "000000000000000000000000",
10040 => "000000000000000000000000",
10041 => "000000000000000000000000",
10042 => "000000000000000000000000",
10043 => "000000000000000000000000",
10044 => "000000000000000000000000",
10045 => "000000000000000000000000",
10046 => "000000000000000000000000",
10047 => "000000000000000000000000",
10048 => "000000000000000000000000",
10049 => "000000000000000000000000",
10050 => "000000000000000000000000",
10051 => "000000000000000000000000",
10052 => "000000000000000000000000",
10053 => "000000000000000000000000",
10054 => "000000000000000000000000",
10055 => "000000000000000000000000",
10056 => "000000000000000000000000",
10057 => "000000000000000000000000",
10058 => "000000000000000000000000",
10059 => "000000000000000000000000",
10060 => "000000000000000000000000",
10061 => "000000000000000000000000",
10062 => "000000000000000000000000",
10063 => "000000000000000000000000",
10064 => "000000000000000000000000",
10065 => "000000000000000000000000",
10066 => "000000000000000000000000",
10067 => "000000000000000000000000",
10068 => "000000000000000000000000",
10069 => "000000000000000000000000",
10070 => "000000000000000000000000",
10071 => "000000000000000000000000",
10072 => "000000000000000000000000",
10073 => "000000000000000000000000",
10074 => "000000000000000000000000",
10075 => "000000000000000000000000",
10076 => "000000000000000000000000",
10077 => "000000000000000000000000",
10078 => "000000000000000000000000",
10079 => "000000000000000000000000",
10080 => "000000000000000000000000",
10081 => "000000000000000000000000",
10082 => "000000000000000000000000",
10083 => "000000000000000000000000",
10084 => "000000000000000000000000",
10085 => "000000000000000000000000",
10086 => "000000000000000000000000",
10087 => "000000000000000000000000",
10088 => "000000000000000000000000",
10089 => "000000000000000000000000",
10090 => "000000000000000000000000",
10091 => "000000000000000000000000",
10092 => "000000000000000000000000",
10093 => "000000000000000000000000",
10094 => "000000010000000100000001",
10095 => "000000110000001100000011",
10096 => "000000110000001100000011",
10097 => "000000000000000000000000",
10098 => "000000000000000000000000",
10099 => "000000000000000000000000",
10100 => "000000000000000000000000",
10101 => "000000000000000000000000",
10102 => "000000000000000000000000",
10103 => "000001100000011000000110",
10104 => "010000110100001101000011",
10105 => "010000110100001101000011",
10106 => "010111110101111101011111",
10107 => "011001100110011001100110",
10108 => "001111010011110100111101",
10109 => "000000000000000000000000",
10110 => "000001000000010000000100",
10111 => "010000110100001101000011",
10112 => "010000110100001101000011",
10113 => "010000110100001101000011",
10114 => "010000110100001101000011",
10115 => "010000110100001101000011",
10116 => "010000110100001101000011",
10117 => "010000110100001101000011",
10118 => "010000110100001101000011",
10119 => "010000110100001101000011",
10120 => "010000110100001101000011",
10121 => "010000110100001101000011",
10122 => "010000110100001101000011",
10123 => "010000110100001101000011",
10124 => "010000110100001101000011",
10125 => "010000110100001101000011",
10126 => "010000110100001101000011",
10127 => "000101110001011100010111",
10128 => "000000000000000000000000",
10129 => "001000000010000000100000",
10130 => "011001100110011001100110",
10131 => "011001100110011001100110",
10132 => "010000110100001101000011",
10133 => "010000110100001101000011",
10134 => "000110010001100100011001",
10135 => "000000000000000000000000",
10136 => "000000000000000000000000",
10137 => "000000000000000000000000",
10138 => "000000000000000000000000",
10139 => "000000000000000000000000",
10140 => "000000000000000000000000",
10141 => "000000100000001000000010",
10142 => "000000110000001100000011",
10143 => "000000100000001000000010",
10144 => "000000000000000000000000",
10145 => "000000000000000000000000",
10146 => "000000000000000000000000",
10147 => "000000000000000000000000",
10148 => "000000000000000000000000",
10149 => "000000000000000000000000",
10150 => "000000000000000000000000",
10151 => "000000000000000000000000",
10152 => "000000000000000000000000",
10153 => "000000000000000000000000",
10154 => "000000000000000000000000",
10155 => "000000000000000000000000",
10156 => "000000000000000000000000",
10157 => "000000000000000000000000",
10158 => "000000000000000000000000",
10159 => "000000000000000000000000",
10160 => "000000000000000000000000",
10161 => "000000000000000000000000",
10162 => "000000000000000000000000",
10163 => "000000000000000000000000",
10164 => "000000000000000000000000",
10165 => "000000000000000000000000",
10166 => "000000000000000000000000",
10167 => "000000000000000000000000",
10168 => "000000000000000000000000",
10169 => "000000000000000000000000",
10170 => "000000000000000000000000",
10171 => "000000000000000000000000",
10172 => "000000000000000000000000",
10173 => "000000000000000000000000",
10174 => "000000000000000000000000",
10175 => "000000000000000000000000",
10176 => "000000000000000000000000",
10177 => "000000000000000000000000",
10178 => "000000000000000000000000",
10179 => "000000000000000000000000",
10180 => "000000000000000000000000",
10181 => "000000000000000000000000",
10182 => "000000000000000000000000",
10183 => "000000000000000000000000",
10184 => "000000000000000000000000",
10185 => "000000000000000000000000",
10186 => "000000000000000000000000",
10187 => "000000000000000000000000",
10188 => "000000000000000000000000",
10189 => "000000000000000000000000",
10190 => "000000000000000000000000",
10191 => "000000000000000000000000",
10192 => "000000000000000000000000",
10193 => "000000000000000000000000",
10194 => "000000000000000000000000",
10195 => "000000000000000000000000",
10196 => "000000000000000000000000",
10197 => "000000000000000000000000",
10198 => "000000000000000000000000",
10199 => "000000000000000000000000",
10200 => "000000000000000000000000",
10201 => "000000000000000000000000",
10202 => "000000000000000000000000",
10203 => "000000000000000000000000",
10204 => "000000000000000000000000",
10205 => "000000000000000000000000",
10206 => "000000000000000000000000",
10207 => "000000000000000000000000",
10208 => "000000000000000000000000",
10209 => "000000000000000000000000",
10210 => "000000000000000000000000",
10211 => "000000000000000000000000",
10212 => "000000000000000000000000",
10213 => "000000000000000000000000",
10214 => "000000000000000000000000",
10215 => "000000000000000000000000",
10216 => "000000000000000000000000",
10217 => "000000000000000000000000",
10218 => "000000000000000000000000",
10219 => "000000000000000000000000",
10220 => "000000000000000000000000",
10221 => "000000000000000000000000",
10222 => "000000000000000000000000",
10223 => "000000000000000000000000",
10224 => "000000000000000000000000",
10225 => "000000000000000000000000",
10226 => "000000000000000000000000",
10227 => "000000000000000000000000",
10228 => "000000000000000000000000",
10229 => "000000000000000000000000",
10230 => "000000000000000000000000",
10231 => "000000000000000000000000",
10232 => "000000000000000000000000",
10233 => "000000000000000000000000",
10234 => "000000000000000000000000",
10235 => "000000000000000000000000",
10236 => "000000000000000000000000",
10237 => "000000000000000000000000",
10238 => "000000000000000000000000",
10239 => "000000000000000000000000",
10240 => "000000000000000000000000",
10241 => "000000000000000000000000",
10242 => "000000000000000000000000",
10243 => "000000000000000000000000",
10244 => "001100000011000000110000",
10245 => "011001100110011001100110",
10246 => "010110010101100101011001",
10247 => "000000000000000000000000",
10248 => "000000000000000000000000",
10249 => "000000000000000000000000",
10250 => "000000000000000000000000",
10251 => "000000000000000000000000",
10252 => "000000000000000000000000",
10253 => "000001100000011000000110",
10254 => "010000110100001101000011",
10255 => "010000110100001101000011",
10256 => "010111110101111101011111",
10257 => "011001100110011001100110",
10258 => "001111010011110100111101",
10259 => "000000000000000000000000",
10260 => "000001000000010000000100",
10261 => "010000110100001101000011",
10262 => "010000110100001101000011",
10263 => "010000110100001101000011",
10264 => "010000110100001101000011",
10265 => "010000110100001101000011",
10266 => "010000110100001101000011",
10267 => "010000110100001101000011",
10268 => "010000110100001101000011",
10269 => "010000110100001101000011",
10270 => "010000110100001101000011",
10271 => "010000110100001101000011",
10272 => "010000110100001101000011",
10273 => "010000110100001101000011",
10274 => "010000110100001101000011",
10275 => "010000110100001101000011",
10276 => "010000110100001101000011",
10277 => "000101110001011100010111",
10278 => "000000000000000000000000",
10279 => "001000000010000000100000",
10280 => "011001100110011001100110",
10281 => "011001100110011001100110",
10282 => "010000110100001101000011",
10283 => "010000110100001101000011",
10284 => "000110010001100100011001",
10285 => "000000000000000000000000",
10286 => "000000000000000000000000",
10287 => "000000000000000000000000",
10288 => "000000000000000000000000",
10289 => "000000000000000000000000",
10290 => "000000000000000000000000",
10291 => "001111010011110100111101",
10292 => "011001100110011001100110",
10293 => "010011010100110101001101",
10294 => "000000000000000000000000",
10295 => "000000000000000000000000",
10296 => "000000000000000000000000",
10297 => "000000000000000000000000",
10298 => "000000000000000000000000",
10299 => "000000000000000000000000",
10300 => "000000000000000000000000",
10301 => "000000000000000000000000",
10302 => "000000000000000000000000",
10303 => "000000000000000000000000",
10304 => "000000000000000000000000",
10305 => "000000000000000000000000",
10306 => "000000000000000000000000",
10307 => "000000000000000000000000",
10308 => "000000000000000000000000",
10309 => "000000000000000000000000",
10310 => "000000000000000000000000",
10311 => "000000000000000000000000",
10312 => "000000000000000000000000",
10313 => "000000000000000000000000",
10314 => "000000000000000000000000",
10315 => "000000000000000000000000",
10316 => "000000000000000000000000",
10317 => "000000000000000000000000",
10318 => "000000000000000000000000",
10319 => "000000000000000000000000",
10320 => "000000000000000000000000",
10321 => "000000000000000000000000",
10322 => "000000000000000000000000",
10323 => "000000000000000000000000",
10324 => "000000000000000000000000",
10325 => "000000000000000000000000",
10326 => "000000000000000000000000",
10327 => "000000000000000000000000",
10328 => "000000000000000000000000",
10329 => "000000000000000000000000",
10330 => "000000000000000000000000",
10331 => "000000000000000000000000",
10332 => "000000000000000000000000",
10333 => "000000000000000000000000",
10334 => "000000000000000000000000",
10335 => "000000000000000000000000",
10336 => "000000000000000000000000",
10337 => "000000000000000000000000",
10338 => "000000000000000000000000",
10339 => "000000000000000000000000",
10340 => "000000000000000000000000",
10341 => "000000000000000000000000",
10342 => "000000000000000000000000",
10343 => "000000000000000000000000",
10344 => "000000000000000000000000",
10345 => "000000000000000000000000",
10346 => "000000000000000000000000",
10347 => "000000000000000000000000",
10348 => "000000000000000000000000",
10349 => "000000000000000000000000",
10350 => "000000000000000000000000",
10351 => "000000000000000000000000",
10352 => "000000000000000000000000",
10353 => "000000000000000000000000",
10354 => "000000000000000000000000",
10355 => "000000000000000000000000",
10356 => "000000000000000000000000",
10357 => "000000000000000000000000",
10358 => "000000000000000000000000",
10359 => "000000000000000000000000",
10360 => "000000000000000000000000",
10361 => "000000000000000000000000",
10362 => "000000000000000000000000",
10363 => "000000000000000000000000",
10364 => "000000000000000000000000",
10365 => "000000000000000000000000",
10366 => "000000000000000000000000",
10367 => "000000000000000000000000",
10368 => "000000000000000000000000",
10369 => "000000000000000000000000",
10370 => "000000000000000000000000",
10371 => "000000000000000000000000",
10372 => "000000000000000000000000",
10373 => "000000000000000000000000",
10374 => "000000000000000000000000",
10375 => "000000000000000000000000",
10376 => "000000000000000000000000",
10377 => "000000000000000000000000",
10378 => "000000000000000000000000",
10379 => "000000000000000000000000",
10380 => "000000000000000000000000",
10381 => "000000000000000000000000",
10382 => "000000000000000000000000",
10383 => "000000000000000000000000",
10384 => "000000000000000000000000",
10385 => "000000000000000000000000",
10386 => "000000000000000000000000",
10387 => "000000000000000000000000",
10388 => "000000000000000000000000",
10389 => "000000000000000000000000",
10390 => "000000000000000000000000",
10391 => "000000000000000000000000",
10392 => "000000000000000000000000",
10393 => "000000000000000000000000",
10394 => "001100000011000000110000",
10395 => "011001100110011001100110",
10396 => "010110010101100101011001",
10397 => "000000000000000000000000",
10398 => "000000000000000000000000",
10399 => "000000000000000000000000",
10400 => "000000000000000000000000",
10401 => "000000000000000000000000",
10402 => "000000000000000000000000",
10403 => "000001100000011000000110",
10404 => "010000110100001101000011",
10405 => "010000110100001101000011",
10406 => "010111110101111101011111",
10407 => "011001100110011001100110",
10408 => "001111010011110100111101",
10409 => "000000000000000000000000",
10410 => "000001000000010000000100",
10411 => "010000110100001101000011",
10412 => "010000110100001101000011",
10413 => "010000110100001101000011",
10414 => "010000110100001101000011",
10415 => "010000110100001101000011",
10416 => "010000110100001101000011",
10417 => "010000110100001101000011",
10418 => "010000110100001101000011",
10419 => "010000110100001101000011",
10420 => "010000110100001101000011",
10421 => "010000110100001101000011",
10422 => "010000110100001101000011",
10423 => "010000110100001101000011",
10424 => "010000110100001101000011",
10425 => "010000110100001101000011",
10426 => "010000110100001101000011",
10427 => "000101110001011100010111",
10428 => "000000000000000000000000",
10429 => "001000000010000000100000",
10430 => "011001100110011001100110",
10431 => "011001100110011001100110",
10432 => "010000110100001101000011",
10433 => "010000110100001101000011",
10434 => "000110010001100100011001",
10435 => "000000000000000000000000",
10436 => "000000000000000000000000",
10437 => "000000000000000000000000",
10438 => "000000000000000000000000",
10439 => "000000000000000000000000",
10440 => "000000000000000000000000",
10441 => "001111010011110100111101",
10442 => "011001100110011001100110",
10443 => "010011010100110101001101",
10444 => "000000000000000000000000",
10445 => "000000000000000000000000",
10446 => "000000000000000000000000",
10447 => "000000000000000000000000",
10448 => "000000000000000000000000",
10449 => "000000000000000000000000",
10450 => "000000000000000000000000",
10451 => "000000000000000000000000",
10452 => "000000000000000000000000",
10453 => "000000000000000000000000",
10454 => "000000000000000000000000",
10455 => "000000000000000000000000",
10456 => "000000000000000000000000",
10457 => "000000000000000000000000",
10458 => "000000000000000000000000",
10459 => "000000000000000000000000",
10460 => "000000000000000000000000",
10461 => "000000000000000000000000",
10462 => "000000000000000000000000",
10463 => "000000000000000000000000",
10464 => "000000000000000000000000",
10465 => "000000000000000000000000",
10466 => "000000000000000000000000",
10467 => "000000000000000000000000",
10468 => "000000000000000000000000",
10469 => "000000000000000000000000",
10470 => "000000000000000000000000",
10471 => "000000000000000000000000",
10472 => "000000000000000000000000",
10473 => "000000000000000000000000",
10474 => "000000000000000000000000",
10475 => "000000000000000000000000",
10476 => "000000000000000000000000",
10477 => "000000000000000000000000",
10478 => "000000000000000000000000",
10479 => "000000000000000000000000",
10480 => "000000000000000000000000",
10481 => "000000000000000000000000",
10482 => "000000000000000000000000",
10483 => "000000000000000000000000",
10484 => "000000000000000000000000",
10485 => "000000000000000000000000",
10486 => "000000000000000000000000",
10487 => "000000000000000000000000",
10488 => "000000000000000000000000",
10489 => "000000000000000000000000",
10490 => "000000000000000000000000",
10491 => "000000000000000000000000",
10492 => "000000000000000000000000",
10493 => "000000000000000000000000",
10494 => "000000000000000000000000",
10495 => "000000000000000000000000",
10496 => "000000000000000000000000",
10497 => "000000000000000000000000",
10498 => "000000000000000000000000",
10499 => "000000000000000000000000",
10500 => "000000000000000000000000",
10501 => "000000000000000000000000",
10502 => "000000000000000000000000",
10503 => "000000000000000000000000",
10504 => "000000000000000000000000",
10505 => "000000000000000000000000",
10506 => "000000000000000000000000",
10507 => "000000000000000000000000",
10508 => "000000000000000000000000",
10509 => "000000000000000000000000",
10510 => "000000000000000000000000",
10511 => "000000000000000000000000",
10512 => "000000000000000000000000",
10513 => "000000000000000000000000",
10514 => "000000000000000000000000",
10515 => "000000000000000000000000",
10516 => "000000000000000000000000",
10517 => "000000000000000000000000",
10518 => "000000000000000000000000",
10519 => "000000000000000000000000",
10520 => "000000000000000000000000",
10521 => "000000000000000000000000",
10522 => "000000000000000000000000",
10523 => "000000000000000000000000",
10524 => "000000000000000000000000",
10525 => "000000000000000000000000",
10526 => "000000000000000000000000",
10527 => "000000000000000000000000",
10528 => "000000000000000000000000",
10529 => "000000000000000000000000",
10530 => "000000000000000000000000",
10531 => "000000000000000000000000",
10532 => "000000000000000000000000",
10533 => "000000000000000000000000",
10534 => "000000000000000000000000",
10535 => "000000000000000000000000",
10536 => "000000000000000000000000",
10537 => "000000000000000000000000",
10538 => "000000000000000000000000",
10539 => "000000000000000000000000",
10540 => "000000000000000000000000",
10541 => "000000000000000000000000",
10542 => "000000000000000000000000",
10543 => "000000000000000000000000",
10544 => "001100000011000000110000",
10545 => "011001100110011001100110",
10546 => "010110010101100101011001",
10547 => "000000000000000000000000",
10548 => "000000000000000000000000",
10549 => "000000000000000000000000",
10550 => "000000000000000000000000",
10551 => "000000000000000000000000",
10552 => "000000000000000000000000",
10553 => "000001100000011000000110",
10554 => "010000110100001101000011",
10555 => "010000110100001101000011",
10556 => "010111110101111101011111",
10557 => "011001100110011001100110",
10558 => "010011110100111101001111",
10559 => "001011100010111000101110",
10560 => "001011110010111100101111",
10561 => "010000110100001101000011",
10562 => "010000110100001101000011",
10563 => "010000110100001101000011",
10564 => "010000110100001101000011",
10565 => "010000110100001101000011",
10566 => "010000110100001101000011",
10567 => "010000110100001101000011",
10568 => "010000110100001101000011",
10569 => "010000110100001101000011",
10570 => "010000110100001101000011",
10571 => "010000110100001101000011",
10572 => "010000110100001101000011",
10573 => "010000110100001101000011",
10574 => "010000110100001101000011",
10575 => "010000110100001101000011",
10576 => "010000110100001101000011",
10577 => "001101010011010100110101",
10578 => "001011100010111000101110",
10579 => "010000000100000001000000",
10580 => "011001100110011001100110",
10581 => "011001100110011001100110",
10582 => "010000110100001101000011",
10583 => "010000110100001101000011",
10584 => "000110010001100100011001",
10585 => "000000000000000000000000",
10586 => "000000000000000000000000",
10587 => "000000000000000000000000",
10588 => "000000000000000000000000",
10589 => "000000000000000000000000",
10590 => "000000000000000000000000",
10591 => "001111010011110100111101",
10592 => "011001100110011001100110",
10593 => "010011010100110101001101",
10594 => "000000000000000000000000",
10595 => "000000000000000000000000",
10596 => "000000000000000000000000",
10597 => "000000000000000000000000",
10598 => "000000000000000000000000",
10599 => "000000000000000000000000",
10600 => "000000000000000000000000",
10601 => "000000000000000000000000",
10602 => "000000000000000000000000",
10603 => "000000000000000000000000",
10604 => "000000000000000000000000",
10605 => "000000000000000000000000",
10606 => "000000000000000000000000",
10607 => "000000000000000000000000",
10608 => "000000000000000000000000",
10609 => "000000000000000000000000",
10610 => "000000000000000000000000",
10611 => "000000000000000000000000",
10612 => "000000000000000000000000",
10613 => "000000000000000000000000",
10614 => "000000000000000000000000",
10615 => "000000000000000000000000",
10616 => "000000000000000000000000",
10617 => "000000000000000000000000",
10618 => "000000000000000000000000",
10619 => "000000000000000000000000",
10620 => "000000000000000000000000",
10621 => "000000000000000000000000",
10622 => "000000000000000000000000",
10623 => "000000000000000000000000",
10624 => "000000000000000000000000",
10625 => "000000000000000000000000",
10626 => "000000000000000000000000",
10627 => "000000000000000000000000",
10628 => "000000000000000000000000",
10629 => "000000000000000000000000",
10630 => "000000000000000000000000",
10631 => "000000000000000000000000",
10632 => "000000000000000000000000",
10633 => "000000000000000000000000",
10634 => "000000000000000000000000",
10635 => "000000000000000000000000",
10636 => "000000000000000000000000",
10637 => "000000000000000000000000",
10638 => "000000000000000000000000",
10639 => "000000000000000000000000",
10640 => "000000000000000000000000",
10641 => "000000000000000000000000",
10642 => "000000000000000000000000",
10643 => "000000000000000000000000",
10644 => "000000000000000000000000",
10645 => "000000000000000000000000",
10646 => "000000000000000000000000",
10647 => "000000000000000000000000",
10648 => "000000000000000000000000",
10649 => "000000000000000000000000",
10650 => "000000000000000000000000",
10651 => "000000000000000000000000",
10652 => "000000000000000000000000",
10653 => "000000000000000000000000",
10654 => "000000000000000000000000",
10655 => "000000000000000000000000",
10656 => "000000000000000000000000",
10657 => "000000000000000000000000",
10658 => "000000000000000000000000",
10659 => "000000000000000000000000",
10660 => "000000000000000000000000",
10661 => "000000000000000000000000",
10662 => "000000000000000000000000",
10663 => "000000000000000000000000",
10664 => "000000000000000000000000",
10665 => "000000000000000000000000",
10666 => "000000000000000000000000",
10667 => "000000000000000000000000",
10668 => "000000000000000000000000",
10669 => "000000000000000000000000",
10670 => "000000000000000000000000",
10671 => "000000000000000000000000",
10672 => "000000000000000000000000",
10673 => "000000000000000000000000",
10674 => "000000000000000000000000",
10675 => "000000000000000000000000",
10676 => "000000000000000000000000",
10677 => "000000000000000000000000",
10678 => "000000000000000000000000",
10679 => "000000000000000000000000",
10680 => "000000000000000000000000",
10681 => "000000000000000000000000",
10682 => "000000000000000000000000",
10683 => "000000000000000000000000",
10684 => "000000000000000000000000",
10685 => "000000000000000000000000",
10686 => "000000000000000000000000",
10687 => "000000000000000000000000",
10688 => "000000000000000000000000",
10689 => "000000000000000000000000",
10690 => "000000000000000000000000",
10691 => "000000000000000000000000",
10692 => "000000000000000000000000",
10693 => "000000000000000000000000",
10694 => "001100000011000000110000",
10695 => "011001100110011001100110",
10696 => "010110010101100101011001",
10697 => "000000000000000000000000",
10698 => "000000000000000000000000",
10699 => "000000000000000000000000",
10700 => "000000000000000000000000",
10701 => "000000000000000000000000",
10702 => "000000000000000000000000",
10703 => "000001100000011000000110",
10704 => "010000110100001101000011",
10705 => "010000110100001101000011",
10706 => "010111110101111101011111",
10707 => "011001100110011001100110",
10708 => "010110000101100001011000",
10709 => "010000110100001101000011",
10710 => "010000110100001101000011",
10711 => "010000110100001101000011",
10712 => "010000110100001101000011",
10713 => "010000110100001101000011",
10714 => "010000110100001101000011",
10715 => "010000110100001101000011",
10716 => "010000110100001101000011",
10717 => "010000110100001101000011",
10718 => "010000110100001101000011",
10719 => "010000110100001101000011",
10720 => "010000110100001101000011",
10721 => "010000110100001101000011",
10722 => "010000110100001101000011",
10723 => "010000110100001101000011",
10724 => "010000110100001101000011",
10725 => "010000110100001101000011",
10726 => "010000110100001101000011",
10727 => "010000110100001101000011",
10728 => "010000110100001101000011",
10729 => "010011100100111001001110",
10730 => "011001100110011001100110",
10731 => "011001100110011001100110",
10732 => "010000110100001101000011",
10733 => "010000110100001101000011",
10734 => "000110010001100100011001",
10735 => "000000000000000000000000",
10736 => "000000000000000000000000",
10737 => "000000000000000000000000",
10738 => "000000000000000000000000",
10739 => "000000000000000000000000",
10740 => "000000000000000000000000",
10741 => "001111010011110100111101",
10742 => "011001100110011001100110",
10743 => "010011010100110101001101",
10744 => "000000000000000000000000",
10745 => "000000000000000000000000",
10746 => "000000000000000000000000",
10747 => "000000000000000000000000",
10748 => "000000000000000000000000",
10749 => "000000000000000000000000",
10750 => "000000000000000000000000",
10751 => "000000000000000000000000",
10752 => "000000000000000000000000",
10753 => "000000000000000000000000",
10754 => "000000000000000000000000",
10755 => "000000000000000000000000",
10756 => "000000000000000000000000",
10757 => "000000000000000000000000",
10758 => "000000000000000000000000",
10759 => "000000000000000000000000",
10760 => "000000000000000000000000",
10761 => "000000000000000000000000",
10762 => "000000000000000000000000",
10763 => "000000000000000000000000",
10764 => "000000000000000000000000",
10765 => "000000000000000000000000",
10766 => "000000000000000000000000",
10767 => "000000000000000000000000",
10768 => "000000000000000000000000",
10769 => "000000000000000000000000",
10770 => "000000000000000000000000",
10771 => "000000000000000000000000",
10772 => "000000000000000000000000",
10773 => "000000000000000000000000",
10774 => "000000000000000000000000",
10775 => "000000000000000000000000",
10776 => "000000000000000000000000",
10777 => "000000000000000000000000",
10778 => "000000000000000000000000",
10779 => "000000000000000000000000",
10780 => "000000000000000000000000",
10781 => "000000000000000000000000",
10782 => "000000000000000000000000",
10783 => "000000000000000000000000",
10784 => "000000000000000000000000",
10785 => "000000000000000000000000",
10786 => "000000000000000000000000",
10787 => "000000000000000000000000",
10788 => "000000000000000000000000",
10789 => "000000000000000000000000",
10790 => "000000000000000000000000",
10791 => "000000000000000000000000",
10792 => "000000000000000000000000",
10793 => "000000000000000000000000",
10794 => "000000000000000000000000",
10795 => "000000000000000000000000",
10796 => "000000000000000000000000",
10797 => "000000000000000000000000",
10798 => "000000000000000000000000",
10799 => "000000000000000000000000",
10800 => "000000000000000000000000",
10801 => "000000000000000000000000",
10802 => "000000000000000000000000",
10803 => "000000000000000000000000",
10804 => "000000000000000000000000",
10805 => "000000000000000000000000",
10806 => "000000000000000000000000",
10807 => "000000000000000000000000",
10808 => "000000000000000000000000",
10809 => "000000000000000000000000",
10810 => "000000000000000000000000",
10811 => "000000000000000000000000",
10812 => "000000000000000000000000",
10813 => "000000000000000000000000",
10814 => "000000000000000000000000",
10815 => "000000000000000000000000",
10816 => "000000000000000000000000",
10817 => "000000000000000000000000",
10818 => "000000000000000000000000",
10819 => "000000000000000000000000",
10820 => "000000000000000000000000",
10821 => "000000000000000000000000",
10822 => "000000000000000000000000",
10823 => "000000000000000000000000",
10824 => "000000000000000000000000",
10825 => "000000000000000000000000",
10826 => "000000000000000000000000",
10827 => "000000000000000000000000",
10828 => "000000000000000000000000",
10829 => "000000000000000000000000",
10830 => "000000000000000000000000",
10831 => "000000000000000000000000",
10832 => "000000000000000000000000",
10833 => "000000000000000000000000",
10834 => "000000000000000000000000",
10835 => "000000000000000000000000",
10836 => "000000000000000000000000",
10837 => "000000000000000000000000",
10838 => "000000000000000000000000",
10839 => "000000000000000000000000",
10840 => "000000000000000000000000",
10841 => "000000000000000000000000",
10842 => "000000000000000000000000",
10843 => "000000000000000000000000",
10844 => "001100000011000000110000",
10845 => "011001100110011001100110",
10846 => "010110010101100101011001",
10847 => "000000000000000000000000",
10848 => "000000000000000000000000",
10849 => "000000000000000000000000",
10850 => "000000000000000000000000",
10851 => "000010100000101000001010",
10852 => "000101110001011100010111",
10853 => "000110110001101100011011",
10854 => "010000110100001101000011",
10855 => "010000110100001101000011",
10856 => "010111110101111101011111",
10857 => "011001100110011001100110",
10858 => "010110000101100001011000",
10859 => "010000110100001101000011",
10860 => "010000110100001101000011",
10861 => "010000110100001101000011",
10862 => "010000110100001101000011",
10863 => "010000110100001101000011",
10864 => "010000110100001101000011",
10865 => "010000110100001101000011",
10866 => "010000110100001101000011",
10867 => "010000110100001101000011",
10868 => "010000110100001101000011",
10869 => "010000110100001101000011",
10870 => "010000110100001101000011",
10871 => "010000110100001101000011",
10872 => "010000110100001101000011",
10873 => "010000110100001101000011",
10874 => "010000110100001101000011",
10875 => "010000110100001101000011",
10876 => "010000110100001101000011",
10877 => "010000110100001101000011",
10878 => "010000110100001101000011",
10879 => "010011100100111001001110",
10880 => "011001100110011001100110",
10881 => "011001100110011001100110",
10882 => "010000110100001101000011",
10883 => "010000110100001101000011",
10884 => "001010000010100000101000",
10885 => "000101110001011100010111",
10886 => "000100010001000100010001",
10887 => "000000000000000000000000",
10888 => "000000000000000000000000",
10889 => "000000000000000000000000",
10890 => "000000000000000000000000",
10891 => "001111010011110100111101",
10892 => "011001100110011001100110",
10893 => "010011010100110101001101",
10894 => "000000000000000000000000",
10895 => "000000000000000000000000",
10896 => "000000000000000000000000",
10897 => "000000000000000000000000",
10898 => "000000000000000000000000",
10899 => "000000000000000000000000",
10900 => "000000000000000000000000",
10901 => "000000000000000000000000",
10902 => "000000000000000000000000",
10903 => "000000000000000000000000",
10904 => "000000000000000000000000",
10905 => "000000000000000000000000",
10906 => "000000000000000000000000",
10907 => "000000000000000000000000",
10908 => "000000000000000000000000",
10909 => "000000000000000000000000",
10910 => "000000000000000000000000",
10911 => "000000000000000000000000",
10912 => "000000000000000000000000",
10913 => "000000000000000000000000",
10914 => "000000000000000000000000",
10915 => "000000000000000000000000",
10916 => "000000000000000000000000",
10917 => "000000000000000000000000",
10918 => "000000000000000000000000",
10919 => "000000000000000000000000",
10920 => "000000000000000000000000",
10921 => "000000000000000000000000",
10922 => "000000000000000000000000",
10923 => "000000000000000000000000",
10924 => "000000000000000000000000",
10925 => "000000000000000000000000",
10926 => "000000000000000000000000",
10927 => "000000000000000000000000",
10928 => "000000000000000000000000",
10929 => "000000000000000000000000",
10930 => "000000000000000000000000",
10931 => "000000000000000000000000",
10932 => "000000000000000000000000",
10933 => "000000000000000000000000",
10934 => "000000000000000000000000",
10935 => "000000000000000000000000",
10936 => "000000000000000000000000",
10937 => "000000000000000000000000",
10938 => "000000000000000000000000",
10939 => "000000000000000000000000",
10940 => "000000000000000000000000",
10941 => "000000000000000000000000",
10942 => "000000000000000000000000",
10943 => "000000000000000000000000",
10944 => "000000000000000000000000",
10945 => "000000000000000000000000",
10946 => "000000000000000000000000",
10947 => "000000000000000000000000",
10948 => "000000000000000000000000",
10949 => "000000000000000000000000",
10950 => "000000000000000000000000",
10951 => "000000000000000000000000",
10952 => "000000000000000000000000",
10953 => "000000000000000000000000",
10954 => "000000000000000000000000",
10955 => "000000000000000000000000",
10956 => "000000000000000000000000",
10957 => "000000000000000000000000",
10958 => "000000000000000000000000",
10959 => "000000000000000000000000",
10960 => "000000000000000000000000",
10961 => "000000000000000000000000",
10962 => "000000000000000000000000",
10963 => "000000000000000000000000",
10964 => "000000000000000000000000",
10965 => "000000000000000000000000",
10966 => "000000000000000000000000",
10967 => "000000000000000000000000",
10968 => "000000000000000000000000",
10969 => "000000000000000000000000",
10970 => "000000000000000000000000",
10971 => "000000000000000000000000",
10972 => "000000000000000000000000",
10973 => "000000000000000000000000",
10974 => "000000000000000000000000",
10975 => "000000000000000000000000",
10976 => "000000000000000000000000",
10977 => "000000000000000000000000",
10978 => "000000000000000000000000",
10979 => "000000000000000000000000",
10980 => "000000000000000000000000",
10981 => "000000000000000000000000",
10982 => "000000000000000000000000",
10983 => "000000000000000000000000",
10984 => "000000000000000000000000",
10985 => "000000000000000000000000",
10986 => "000000000000000000000000",
10987 => "000000000000000000000000",
10988 => "000000000000000000000000",
10989 => "000000000000000000000000",
10990 => "000000000000000000000000",
10991 => "000000000000000000000000",
10992 => "000000000000000000000000",
10993 => "000000000000000000000000",
10994 => "001100000011000000110000",
10995 => "011001100110011001100110",
10996 => "010110010101100101011001",
10997 => "000000000000000000000000",
10998 => "000000000000000000000000",
10999 => "000000000000000000000000",
11000 => "000000000000000000000000",
11001 => "000111010001110100011101",
11002 => "010000110100001101000011",
11003 => "010000110100001101000011",
11004 => "010000110100001101000011",
11005 => "010000110100001101000011",
11006 => "010111110101111101011111",
11007 => "011001100110011001100110",
11008 => "010110000101100001011000",
11009 => "010000110100001101000011",
11010 => "010000110100001101000011",
11011 => "010000110100001101000011",
11012 => "010000110100001101000011",
11013 => "010000110100001101000011",
11014 => "010000110100001101000011",
11015 => "010000110100001101000011",
11016 => "010000110100001101000011",
11017 => "010000110100001101000011",
11018 => "010000110100001101000011",
11019 => "010000110100001101000011",
11020 => "010000110100001101000011",
11021 => "010000110100001101000011",
11022 => "010000110100001101000011",
11023 => "010000110100001101000011",
11024 => "010000110100001101000011",
11025 => "010000110100001101000011",
11026 => "010000110100001101000011",
11027 => "010000110100001101000011",
11028 => "010000110100001101000011",
11029 => "010011100100111001001110",
11030 => "011001100110011001100110",
11031 => "011001100110011001100110",
11032 => "010000110100001101000011",
11033 => "010000110100001101000011",
11034 => "010000110100001101000011",
11035 => "010000110100001101000011",
11036 => "001100000011000000110000",
11037 => "000000000000000000000000",
11038 => "000000000000000000000000",
11039 => "000000000000000000000000",
11040 => "000000000000000000000000",
11041 => "001111010011110100111101",
11042 => "011001100110011001100110",
11043 => "010011010100110101001101",
11044 => "000000000000000000000000",
11045 => "000000000000000000000000",
11046 => "000000000000000000000000",
11047 => "000000000000000000000000",
11048 => "000000000000000000000000",
11049 => "000000000000000000000000",
11050 => "000000000000000000000000",
11051 => "000000000000000000000000",
11052 => "000000000000000000000000",
11053 => "000000000000000000000000",
11054 => "000000000000000000000000",
11055 => "000000000000000000000000",
11056 => "000000000000000000000000",
11057 => "000000000000000000000000",
11058 => "000000000000000000000000",
11059 => "000000000000000000000000",
11060 => "000000000000000000000000",
11061 => "000000000000000000000000",
11062 => "000000000000000000000000",
11063 => "000000000000000000000000",
11064 => "000000000000000000000000",
11065 => "000000000000000000000000",
11066 => "000000000000000000000000",
11067 => "000000000000000000000000",
11068 => "000000000000000000000000",
11069 => "000000000000000000000000",
11070 => "000000000000000000000000",
11071 => "000000000000000000000000",
11072 => "000000000000000000000000",
11073 => "000000000000000000000000",
11074 => "000000000000000000000000",
11075 => "000000000000000000000000",
11076 => "000000000000000000000000",
11077 => "000000000000000000000000",
11078 => "000000000000000000000000",
11079 => "000000000000000000000000",
11080 => "000000000000000000000000",
11081 => "000000000000000000000000",
11082 => "000000000000000000000000",
11083 => "000000000000000000000000",
11084 => "000000000000000000000000",
11085 => "000000000000000000000000",
11086 => "000000000000000000000000",
11087 => "000000000000000000000000",
11088 => "000000000000000000000000",
11089 => "000000000000000000000000",
11090 => "000000000000000000000000",
11091 => "000000000000000000000000",
11092 => "000000000000000000000000",
11093 => "000000000000000000000000",
11094 => "000000000000000000000000",
11095 => "000000000000000000000000",
11096 => "000000000000000000000000",
11097 => "000000000000000000000000",
11098 => "000000000000000000000000",
11099 => "000000000000000000000000",
11100 => "000000000000000000000000",
11101 => "000000000000000000000000",
11102 => "000000000000000000000000",
11103 => "000000000000000000000000",
11104 => "000000000000000000000000",
11105 => "000000000000000000000000",
11106 => "000000000000000000000000",
11107 => "000000000000000000000000",
11108 => "000000000000000000000000",
11109 => "000000000000000000000000",
11110 => "000000000000000000000000",
11111 => "000000000000000000000000",
11112 => "000000000000000000000000",
11113 => "000000000000000000000000",
11114 => "000000000000000000000000",
11115 => "000000000000000000000000",
11116 => "000000000000000000000000",
11117 => "000000000000000000000000",
11118 => "000000000000000000000000",
11119 => "000000000000000000000000",
11120 => "000000000000000000000000",
11121 => "000000000000000000000000",
11122 => "000000000000000000000000",
11123 => "000000000000000000000000",
11124 => "000000000000000000000000",
11125 => "000000000000000000000000",
11126 => "000000000000000000000000",
11127 => "000000000000000000000000",
11128 => "000000000000000000000000",
11129 => "000000000000000000000000",
11130 => "000000000000000000000000",
11131 => "000000000000000000000000",
11132 => "000000000000000000000000",
11133 => "000000000000000000000000",
11134 => "000000000000000000000000",
11135 => "000000000000000000000000",
11136 => "000000000000000000000000",
11137 => "000000000000000000000000",
11138 => "000000000000000000000000",
11139 => "000000000000000000000000",
11140 => "000000000000000000000000",
11141 => "000000000000000000000000",
11142 => "000000000000000000000000",
11143 => "000000000000000000000000",
11144 => "001100000011000000110000",
11145 => "011001100110011001100110",
11146 => "010110010101100101011001",
11147 => "000000000000000000000000",
11148 => "000000000000000000000000",
11149 => "000000000000000000000000",
11150 => "000000000000000000000000",
11151 => "000111010001110100011101",
11152 => "010000110100001101000011",
11153 => "010000110100001101000011",
11154 => "010000110100001101000011",
11155 => "010000110100001101000011",
11156 => "010111110101111101011111",
11157 => "011001100110011001100110",
11158 => "010110000101100001011000",
11159 => "010000110100001101000011",
11160 => "010000110100001101000011",
11161 => "010000110100001101000011",
11162 => "010000110100001101000011",
11163 => "010000110100001101000011",
11164 => "010000110100001101000011",
11165 => "010000110100001101000011",
11166 => "010000110100001101000011",
11167 => "010000110100001101000011",
11168 => "010000110100001101000011",
11169 => "010000110100001101000011",
11170 => "010000110100001101000011",
11171 => "010000110100001101000011",
11172 => "010000110100001101000011",
11173 => "010000110100001101000011",
11174 => "010000110100001101000011",
11175 => "010000110100001101000011",
11176 => "010000110100001101000011",
11177 => "010000110100001101000011",
11178 => "010000110100001101000011",
11179 => "010011100100111001001110",
11180 => "011001100110011001100110",
11181 => "011001100110011001100110",
11182 => "010000110100001101000011",
11183 => "010000110100001101000011",
11184 => "010000110100001101000011",
11185 => "010000110100001101000011",
11186 => "001100000011000000110000",
11187 => "000000000000000000000000",
11188 => "000000000000000000000000",
11189 => "000000000000000000000000",
11190 => "000000000000000000000000",
11191 => "001111010011110100111101",
11192 => "011001100110011001100110",
11193 => "010011010100110101001101",
11194 => "000000000000000000000000",
11195 => "000000000000000000000000",
11196 => "000000000000000000000000",
11197 => "000000000000000000000000",
11198 => "000000000000000000000000",
11199 => "000000000000000000000000",
11200 => "000000000000000000000000",
11201 => "000000000000000000000000",
11202 => "000000000000000000000000",
11203 => "000000000000000000000000",
11204 => "000000000000000000000000",
11205 => "000000000000000000000000",
11206 => "000000000000000000000000",
11207 => "000000000000000000000000",
11208 => "000000000000000000000000",
11209 => "000000000000000000000000",
11210 => "000000000000000000000000",
11211 => "000000000000000000000000",
11212 => "000000000000000000000000",
11213 => "000000000000000000000000",
11214 => "000000000000000000000000",
11215 => "000000000000000000000000",
11216 => "000000000000000000000000",
11217 => "000000000000000000000000",
11218 => "000000000000000000000000",
11219 => "000000000000000000000000",
11220 => "000000000000000000000000",
11221 => "000000000000000000000000",
11222 => "000000000000000000000000",
11223 => "000000000000000000000000",
11224 => "000000000000000000000000",
11225 => "000000000000000000000000",
11226 => "000000000000000000000000",
11227 => "000000000000000000000000",
11228 => "000000000000000000000000",
11229 => "000000000000000000000000",
11230 => "000000000000000000000000",
11231 => "000000000000000000000000",
11232 => "000000000000000000000000",
11233 => "000000000000000000000000",
11234 => "000000000000000000000000",
11235 => "000000000000000000000000",
11236 => "000000000000000000000000",
11237 => "000000000000000000000000",
11238 => "000000000000000000000000",
11239 => "000000000000000000000000",
11240 => "000000000000000000000000",
11241 => "000000000000000000000000",
11242 => "000000000000000000000000",
11243 => "000000000000000000000000",
11244 => "000000000000000000000000",
11245 => "000000000000000000000000",
11246 => "000000000000000000000000",
11247 => "000000000000000000000000",
11248 => "000000000000000000000000",
11249 => "000000000000000000000000",
11250 => "000000000000000000000000",
11251 => "000000000000000000000000",
11252 => "000000000000000000000000",
11253 => "000000000000000000000000",
11254 => "000000000000000000000000",
11255 => "000000000000000000000000",
11256 => "000000000000000000000000",
11257 => "000000000000000000000000",
11258 => "000000000000000000000000",
11259 => "000000000000000000000000",
11260 => "000000000000000000000000",
11261 => "000000000000000000000000",
11262 => "000000000000000000000000",
11263 => "000000000000000000000000",
11264 => "000000000000000000000000",
11265 => "000000000000000000000000",
11266 => "000000000000000000000000",
11267 => "000000000000000000000000",
11268 => "000000000000000000000000",
11269 => "000000000000000000000000",
11270 => "000000000000000000000000",
11271 => "000000000000000000000000",
11272 => "000000000000000000000000",
11273 => "000000000000000000000000",
11274 => "000000000000000000000000",
11275 => "000000000000000000000000",
11276 => "000000000000000000000000",
11277 => "000000000000000000000000",
11278 => "000000000000000000000000",
11279 => "000000000000000000000000",
11280 => "000000000000000000000000",
11281 => "000000000000000000000000",
11282 => "000000000000000000000000",
11283 => "000000000000000000000000",
11284 => "000000000000000000000000",
11285 => "000000000000000000000000",
11286 => "000000000000000000000000",
11287 => "000000000000000000000000",
11288 => "000000000000000000000000",
11289 => "000000000000000000000000",
11290 => "000000000000000000000000",
11291 => "000000000000000000000000",
11292 => "000000000000000000000000",
11293 => "000000000000000000000000",
11294 => "001100000011000000110000",
11295 => "011001100110011001100110",
11296 => "010110010101100101011001",
11297 => "000000000000000000000000",
11298 => "000000000000000000000000",
11299 => "001110000011100000111000",
11300 => "010000110100001101000011",
11301 => "010000110100001101000011",
11302 => "010000110100001101000011",
11303 => "010000110100001101000011",
11304 => "010000110100001101000011",
11305 => "010000110100001101000011",
11306 => "010111110101111101011111",
11307 => "011001100110011001100110",
11308 => "010110000101100001011000",
11309 => "010000110100001101000011",
11310 => "010000110100001101000011",
11311 => "010000110100001101000011",
11312 => "010000110100001101000011",
11313 => "010000110100001101000011",
11314 => "010000110100001101000011",
11315 => "010000110100001101000011",
11316 => "010000110100001101000011",
11317 => "010000110100001101000011",
11318 => "010000110100001101000011",
11319 => "010000110100001101000011",
11320 => "010000110100001101000011",
11321 => "010000110100001101000011",
11322 => "010000110100001101000011",
11323 => "010000110100001101000011",
11324 => "010000110100001101000011",
11325 => "010000110100001101000011",
11326 => "010000110100001101000011",
11327 => "010000110100001101000011",
11328 => "010000110100001101000011",
11329 => "010011100100111001001110",
11330 => "011001100110011001100110",
11331 => "011001100110011001100110",
11332 => "010000110100001101000011",
11333 => "010000110100001101000011",
11334 => "010000110100001101000011",
11335 => "010000110100001101000011",
11336 => "010000110100001101000011",
11337 => "010000110100001101000011",
11338 => "010000110100001101000011",
11339 => "000000010000000100000001",
11340 => "000000000000000000000000",
11341 => "001111010011110100111101",
11342 => "011001100110011001100110",
11343 => "010011010100110101001101",
11344 => "000000000000000000000000",
11345 => "000000000000000000000000",
11346 => "000000000000000000000000",
11347 => "000000000000000000000000",
11348 => "000000000000000000000000",
11349 => "000000000000000000000000",
11350 => "000000000000000000000000",
11351 => "000000000000000000000000",
11352 => "000000000000000000000000",
11353 => "000000000000000000000000",
11354 => "000000000000000000000000",
11355 => "000000000000000000000000",
11356 => "000000000000000000000000",
11357 => "000000000000000000000000",
11358 => "000000000000000000000000",
11359 => "000000000000000000000000",
11360 => "000000000000000000000000",
11361 => "000000000000000000000000",
11362 => "000000000000000000000000",
11363 => "000000000000000000000000",
11364 => "000000000000000000000000",
11365 => "000000000000000000000000",
11366 => "000000000000000000000000",
11367 => "000000000000000000000000",
11368 => "000000000000000000000000",
11369 => "000000000000000000000000",
11370 => "000000000000000000000000",
11371 => "000000000000000000000000",
11372 => "000000000000000000000000",
11373 => "000000000000000000000000",
11374 => "000000000000000000000000",
11375 => "000000000000000000000000",
11376 => "000000000000000000000000",
11377 => "000000000000000000000000",
11378 => "000000000000000000000000",
11379 => "000000000000000000000000",
11380 => "000000000000000000000000",
11381 => "000000000000000000000000",
11382 => "000000000000000000000000",
11383 => "000000000000000000000000",
11384 => "000000000000000000000000",
11385 => "000000000000000000000000",
11386 => "000000000000000000000000",
11387 => "000000000000000000000000",
11388 => "000000000000000000000000",
11389 => "000000000000000000000000",
11390 => "000000000000000000000000",
11391 => "000000000000000000000000",
11392 => "000000000000000000000000",
11393 => "000000000000000000000000",
11394 => "000000000000000000000000",
11395 => "000000000000000000000000",
11396 => "000000000000000000000000",
11397 => "000000000000000000000000",
11398 => "000000000000000000000000",
11399 => "000000000000000000000000",
11400 => "000000000000000000000000",
11401 => "000000000000000000000000",
11402 => "000000000000000000000000",
11403 => "000000000000000000000000",
11404 => "000000000000000000000000",
11405 => "000000000000000000000000",
11406 => "000000000000000000000000",
11407 => "000000000000000000000000",
11408 => "000000000000000000000000",
11409 => "000000000000000000000000",
11410 => "000000000000000000000000",
11411 => "000000000000000000000000",
11412 => "000000000000000000000000",
11413 => "000000000000000000000000",
11414 => "000000000000000000000000",
11415 => "000000000000000000000000",
11416 => "000000000000000000000000",
11417 => "000000000000000000000000",
11418 => "000000000000000000000000",
11419 => "000000000000000000000000",
11420 => "000000000000000000000000",
11421 => "000000000000000000000000",
11422 => "000000000000000000000000",
11423 => "000000000000000000000000",
11424 => "000000000000000000000000",
11425 => "000000000000000000000000",
11426 => "000000000000000000000000",
11427 => "000000000000000000000000",
11428 => "000000000000000000000000",
11429 => "000000000000000000000000",
11430 => "000000000000000000000000",
11431 => "000000000000000000000000",
11432 => "000000000000000000000000",
11433 => "000000000000000000000000",
11434 => "000000000000000000000000",
11435 => "000000000000000000000000",
11436 => "000000000000000000000000",
11437 => "000000000000000000000000",
11438 => "000000000000000000000000",
11439 => "000000000000000000000000",
11440 => "000000000000000000000000",
11441 => "000000000000000000000000",
11442 => "000000000000000000000000",
11443 => "000000000000000000000000",
11444 => "001100000011000000110000",
11445 => "011001100110011001100110",
11446 => "010110010101100101011001",
11447 => "000000000000000000000000",
11448 => "000000000000000000000000",
11449 => "001110000011100000111000",
11450 => "010000110100001101000011",
11451 => "010000110100001101000011",
11452 => "010000110100001101000011",
11453 => "010000110100001101000011",
11454 => "010000110100001101000011",
11455 => "010000110100001101000011",
11456 => "010111110101111101011111",
11457 => "011001100110011001100110",
11458 => "010110000101100001011000",
11459 => "010000110100001101000011",
11460 => "010000110100001101000011",
11461 => "010000110100001101000011",
11462 => "010000110100001101000011",
11463 => "010000110100001101000011",
11464 => "010000110100001101000011",
11465 => "010000110100001101000011",
11466 => "010000110100001101000011",
11467 => "010000110100001101000011",
11468 => "010000110100001101000011",
11469 => "010000110100001101000011",
11470 => "010000110100001101000011",
11471 => "010000110100001101000011",
11472 => "010000110100001101000011",
11473 => "010000110100001101000011",
11474 => "010000110100001101000011",
11475 => "010000110100001101000011",
11476 => "010000110100001101000011",
11477 => "010000110100001101000011",
11478 => "010000110100001101000011",
11479 => "010011100100111001001110",
11480 => "011001100110011001100110",
11481 => "011001100110011001100110",
11482 => "010000110100001101000011",
11483 => "010000110100001101000011",
11484 => "010000110100001101000011",
11485 => "010000110100001101000011",
11486 => "010000110100001101000011",
11487 => "010000110100001101000011",
11488 => "010000110100001101000011",
11489 => "000000010000000100000001",
11490 => "000000000000000000000000",
11491 => "001111010011110100111101",
11492 => "011001100110011001100110",
11493 => "010011010100110101001101",
11494 => "000000000000000000000000",
11495 => "000000000000000000000000",
11496 => "000000000000000000000000",
11497 => "000000000000000000000000",
11498 => "000000000000000000000000",
11499 => "000000000000000000000000",
11500 => "000000000000000000000000",
11501 => "000000000000000000000000",
11502 => "000000000000000000000000",
11503 => "000000000000000000000000",
11504 => "000000000000000000000000",
11505 => "000000000000000000000000",
11506 => "000000000000000000000000",
11507 => "000000000000000000000000",
11508 => "000000000000000000000000",
11509 => "000000000000000000000000",
11510 => "000000000000000000000000",
11511 => "000000000000000000000000",
11512 => "000000000000000000000000",
11513 => "000000000000000000000000",
11514 => "000000000000000000000000",
11515 => "000000000000000000000000",
11516 => "000000000000000000000000",
11517 => "000000000000000000000000",
11518 => "000000000000000000000000",
11519 => "000000000000000000000000",
11520 => "000000000000000000000000",
11521 => "000000000000000000000000",
11522 => "000000000000000000000000",
11523 => "000000000000000000000000",
11524 => "000000000000000000000000",
11525 => "000000000000000000000000",
11526 => "000000000000000000000000",
11527 => "000000000000000000000000",
11528 => "000000000000000000000000",
11529 => "000000000000000000000000",
11530 => "000000000000000000000000",
11531 => "000000000000000000000000",
11532 => "000000000000000000000000",
11533 => "000000000000000000000000",
11534 => "000000000000000000000000",
11535 => "000000000000000000000000",
11536 => "000000000000000000000000",
11537 => "000000000000000000000000",
11538 => "000000000000000000000000",
11539 => "000000000000000000000000",
11540 => "000000000000000000000000",
11541 => "000000000000000000000000",
11542 => "000000000000000000000000",
11543 => "000000000000000000000000",
11544 => "000000000000000000000000",
11545 => "000000000000000000000000",
11546 => "000000000000000000000000",
11547 => "000000000000000000000000",
11548 => "000000000000000000000000",
11549 => "000000000000000000000000",
11550 => "000000000000000000000000",
11551 => "000000000000000000000000",
11552 => "000000000000000000000000",
11553 => "000000000000000000000000",
11554 => "000000000000000000000000",
11555 => "000000000000000000000000",
11556 => "000000000000000000000000",
11557 => "000000000000000000000000",
11558 => "000000000000000000000000",
11559 => "000000000000000000000000",
11560 => "000000000000000000000000",
11561 => "000000000000000000000000",
11562 => "000000000000000000000000",
11563 => "000000000000000000000000",
11564 => "000000000000000000000000",
11565 => "000000000000000000000000",
11566 => "000000000000000000000000",
11567 => "000000000000000000000000",
11568 => "000000000000000000000000",
11569 => "000000000000000000000000",
11570 => "000000000000000000000000",
11571 => "000000000000000000000000",
11572 => "000000000000000000000000",
11573 => "000000000000000000000000",
11574 => "000000000000000000000000",
11575 => "000000000000000000000000",
11576 => "000000000000000000000000",
11577 => "000000000000000000000000",
11578 => "000000000000000000000000",
11579 => "000000000000000000000000",
11580 => "000000000000000000000000",
11581 => "000000000000000000000000",
11582 => "000000000000000000000000",
11583 => "000000000000000000000000",
11584 => "000000000000000000000000",
11585 => "000000000000000000000000",
11586 => "000000000000000000000000",
11587 => "000000000000000000000000",
11588 => "000000000000000000000000",
11589 => "000000000000000000000000",
11590 => "000000000000000000000000",
11591 => "000000000000000000000000",
11592 => "000000000000000000000000",
11593 => "000000000000000000000000",
11594 => "000100000001000000010000",
11595 => "001000110010001100100011",
11596 => "001001000010010000100100",
11597 => "001011000010110000101100",
11598 => "001011000010110000101100",
11599 => "001111110011111100111111",
11600 => "010000110100001101000011",
11601 => "010000110100001101000011",
11602 => "010000110100001101000011",
11603 => "010000110100001101000011",
11604 => "010000110100001101000011",
11605 => "010000110100001101000011",
11606 => "010111110101111101011111",
11607 => "011001100110011001100110",
11608 => "010110000101100001011000",
11609 => "010000110100001101000011",
11610 => "010000110100001101000011",
11611 => "010000110100001101000011",
11612 => "010000110100001101000011",
11613 => "010000110100001101000011",
11614 => "010000110100001101000011",
11615 => "010000110100001101000011",
11616 => "010000110100001101000011",
11617 => "010000110100001101000011",
11618 => "010000110100001101000011",
11619 => "010000110100001101000011",
11620 => "010000110100001101000011",
11621 => "010000110100001101000011",
11622 => "010000110100001101000011",
11623 => "010000110100001101000011",
11624 => "010000110100001101000011",
11625 => "010000110100001101000011",
11626 => "010000110100001101000011",
11627 => "010000110100001101000011",
11628 => "010000110100001101000011",
11629 => "010011100100111001001110",
11630 => "011001100110011001100110",
11631 => "011001100110011001100110",
11632 => "010000110100001101000011",
11633 => "010000110100001101000011",
11634 => "010000110100001101000011",
11635 => "010000110100001101000011",
11636 => "010000110100001101000011",
11637 => "010000110100001101000011",
11638 => "010000110100001101000011",
11639 => "001011000010110000101100",
11640 => "001011000010110000101100",
11641 => "001001110010011100100111",
11642 => "001000110010001100100011",
11643 => "000110100001101000011010",
11644 => "000000000000000000000000",
11645 => "000000000000000000000000",
11646 => "000000000000000000000000",
11647 => "000000000000000000000000",
11648 => "000000000000000000000000",
11649 => "000000000000000000000000",
11650 => "000000000000000000000000",
11651 => "000000000000000000000000",
11652 => "000000000000000000000000",
11653 => "000000000000000000000000",
11654 => "000000000000000000000000",
11655 => "000000000000000000000000",
11656 => "000000000000000000000000",
11657 => "000000000000000000000000",
11658 => "000000000000000000000000",
11659 => "000000000000000000000000",
11660 => "000000000000000000000000",
11661 => "000000000000000000000000",
11662 => "000000000000000000000000",
11663 => "000000000000000000000000",
11664 => "000000000000000000000000",
11665 => "000000000000000000000000",
11666 => "000000000000000000000000",
11667 => "000000000000000000000000",
11668 => "000000000000000000000000",
11669 => "000000000000000000000000",
11670 => "000000000000000000000000",
11671 => "000000000000000000000000",
11672 => "000000000000000000000000",
11673 => "000000000000000000000000",
11674 => "000000000000000000000000",
11675 => "000000000000000000000000",
11676 => "000000000000000000000000",
11677 => "000000000000000000000000",
11678 => "000000000000000000000000",
11679 => "000000000000000000000000",
11680 => "000000000000000000000000",
11681 => "000000000000000000000000",
11682 => "000000000000000000000000",
11683 => "000000000000000000000000",
11684 => "000000000000000000000000",
11685 => "000000000000000000000000",
11686 => "000000000000000000000000",
11687 => "000000000000000000000000",
11688 => "000000000000000000000000",
11689 => "000000000000000000000000",
11690 => "000000000000000000000000",
11691 => "000000000000000000000000",
11692 => "000000000000000000000000",
11693 => "000000000000000000000000",
11694 => "000000000000000000000000",
11695 => "000000000000000000000000",
11696 => "000000000000000000000000",
11697 => "000000000000000000000000",
11698 => "000000000000000000000000",
11699 => "000000000000000000000000",
11700 => "000000000000000000000000",
11701 => "000000000000000000000000",
11702 => "000000000000000000000000",
11703 => "000000000000000000000000",
11704 => "000000000000000000000000",
11705 => "000000000000000000000000",
11706 => "000000000000000000000000",
11707 => "000000000000000000000000",
11708 => "000000000000000000000000",
11709 => "000000000000000000000000",
11710 => "000000000000000000000000",
11711 => "000000000000000000000000",
11712 => "000000000000000000000000",
11713 => "000000000000000000000000",
11714 => "000000000000000000000000",
11715 => "000000000000000000000000",
11716 => "000000000000000000000000",
11717 => "000000000000000000000000",
11718 => "000000000000000000000000",
11719 => "000000000000000000000000",
11720 => "000000000000000000000000",
11721 => "000000000000000000000000",
11722 => "000000000000000000000000",
11723 => "000000000000000000000000",
11724 => "000000000000000000000000",
11725 => "000000000000000000000000",
11726 => "000000000000000000000000",
11727 => "000000000000000000000000",
11728 => "000000000000000000000000",
11729 => "000000000000000000000000",
11730 => "000000000000000000000000",
11731 => "000000000000000000000000",
11732 => "000000000000000000000000",
11733 => "000000000000000000000000",
11734 => "000000000000000000000000",
11735 => "000000000000000000000000",
11736 => "000000000000000000000000",
11737 => "000000000000000000000000",
11738 => "000000000000000000000000",
11739 => "000000000000000000000000",
11740 => "000000000000000000000000",
11741 => "000000000000000000000000",
11742 => "000000000000000000000000",
11743 => "000000000000000000000000",
11744 => "000000000000000000000000",
11745 => "000000000000000000000000",
11746 => "000010000000100000001000",
11747 => "010000110100001101000011",
11748 => "010000110100001101000011",
11749 => "010000110100001101000011",
11750 => "010000110100001101000011",
11751 => "010000110100001101000011",
11752 => "010000110100001101000011",
11753 => "010000110100001101000011",
11754 => "010000110100001101000011",
11755 => "010000110100001101000011",
11756 => "010111110101111101011111",
11757 => "011001100110011001100110",
11758 => "010110000101100001011000",
11759 => "010000110100001101000011",
11760 => "010000110100001101000011",
11761 => "010000110100001101000011",
11762 => "010000110100001101000011",
11763 => "010000110100001101000011",
11764 => "010000110100001101000011",
11765 => "010000110100001101000011",
11766 => "010000110100001101000011",
11767 => "010000110100001101000011",
11768 => "010000110100001101000011",
11769 => "010000110100001101000011",
11770 => "010000110100001101000011",
11771 => "010000110100001101000011",
11772 => "010000110100001101000011",
11773 => "010000110100001101000011",
11774 => "010000110100001101000011",
11775 => "010000110100001101000011",
11776 => "010000110100001101000011",
11777 => "010000110100001101000011",
11778 => "010000110100001101000011",
11779 => "010011100100111001001110",
11780 => "011001100110011001100110",
11781 => "011001100110011001100110",
11782 => "010000110100001101000011",
11783 => "010000110100001101000011",
11784 => "010000110100001101000011",
11785 => "010000110100001101000011",
11786 => "010000110100001101000011",
11787 => "010000110100001101000011",
11788 => "010000110100001101000011",
11789 => "010000110100001101000011",
11790 => "010000110100001101000011",
11791 => "000110110001101100011011",
11792 => "000000000000000000000000",
11793 => "000000000000000000000000",
11794 => "000000000000000000000000",
11795 => "000000000000000000000000",
11796 => "000000000000000000000000",
11797 => "000000000000000000000000",
11798 => "000000000000000000000000",
11799 => "000000000000000000000000",
11800 => "000000000000000000000000",
11801 => "000000000000000000000000",
11802 => "000000000000000000000000",
11803 => "000000000000000000000000",
11804 => "000000000000000000000000",
11805 => "000000000000000000000000",
11806 => "000000000000000000000000",
11807 => "000000000000000000000000",
11808 => "000000000000000000000000",
11809 => "000000000000000000000000",
11810 => "000000000000000000000000",
11811 => "000000000000000000000000",
11812 => "000000000000000000000000",
11813 => "000000000000000000000000",
11814 => "000000000000000000000000",
11815 => "000000000000000000000000",
11816 => "000000000000000000000000",
11817 => "000000000000000000000000",
11818 => "000000000000000000000000",
11819 => "000000000000000000000000",
11820 => "000000000000000000000000",
11821 => "000000000000000000000000",
11822 => "000000000000000000000000",
11823 => "000000000000000000000000",
11824 => "000000000000000000000000",
11825 => "000000000000000000000000",
11826 => "000000000000000000000000",
11827 => "000000000000000000000000",
11828 => "000000000000000000000000",
11829 => "000000000000000000000000",
11830 => "000000000000000000000000",
11831 => "000000000000000000000000",
11832 => "000000000000000000000000",
11833 => "000000000000000000000000",
11834 => "000000000000000000000000",
11835 => "000000000000000000000000",
11836 => "000000000000000000000000",
11837 => "000000000000000000000000",
11838 => "000000000000000000000000",
11839 => "000000000000000000000000",
11840 => "000000000000000000000000",
11841 => "000000000000000000000000",
11842 => "000000000000000000000000",
11843 => "000000000000000000000000",
11844 => "000000000000000000000000",
11845 => "000000000000000000000000",
11846 => "000000000000000000000000",
11847 => "000000000000000000000000",
11848 => "000000000000000000000000",
11849 => "000000000000000000000000",
11850 => "000000000000000000000000",
11851 => "000000000000000000000000",
11852 => "000000000000000000000000",
11853 => "000000000000000000000000",
11854 => "000000000000000000000000",
11855 => "000000000000000000000000",
11856 => "000000000000000000000000",
11857 => "000000000000000000000000",
11858 => "000000000000000000000000",
11859 => "000000000000000000000000",
11860 => "000000000000000000000000",
11861 => "000000000000000000000000",
11862 => "000000000000000000000000",
11863 => "000000000000000000000000",
11864 => "000000000000000000000000",
11865 => "000000000000000000000000",
11866 => "000000000000000000000000",
11867 => "000000000000000000000000",
11868 => "000000000000000000000000",
11869 => "000000000000000000000000",
11870 => "000000000000000000000000",
11871 => "000000000000000000000000",
11872 => "000000000000000000000000",
11873 => "000000000000000000000000",
11874 => "000000000000000000000000",
11875 => "000000000000000000000000",
11876 => "000000000000000000000000",
11877 => "000000000000000000000000",
11878 => "000000000000000000000000",
11879 => "000000000000000000000000",
11880 => "000000000000000000000000",
11881 => "000000000000000000000000",
11882 => "000000000000000000000000",
11883 => "000000000000000000000000",
11884 => "000000000000000000000000",
11885 => "000000000000000000000000",
11886 => "000000000000000000000000",
11887 => "000000000000000000000000",
11888 => "000000000000000000000000",
11889 => "000000000000000000000000",
11890 => "000000000000000000000000",
11891 => "000000000000000000000000",
11892 => "000111000001110000011100",
11893 => "001000000010000000100000",
11894 => "000110110001101100011011",
11895 => "000101010001010100010101",
11896 => "000110110001101100011011",
11897 => "010000110100001101000011",
11898 => "010000110100001101000011",
11899 => "010000110100001101000011",
11900 => "010000110100001101000011",
11901 => "010000110100001101000011",
11902 => "010000110100001101000011",
11903 => "010000110100001101000011",
11904 => "010000110100001101000011",
11905 => "010000110100001101000011",
11906 => "010111110101111101011111",
11907 => "011001100110011001100110",
11908 => "010110000101100001011000",
11909 => "010000110100001101000011",
11910 => "010000110100001101000011",
11911 => "010000110100001101000011",
11912 => "010000110100001101000011",
11913 => "010000110100001101000011",
11914 => "010000110100001101000011",
11915 => "010000110100001101000011",
11916 => "010000110100001101000011",
11917 => "010000110100001101000011",
11918 => "010000110100001101000011",
11919 => "010000110100001101000011",
11920 => "010000110100001101000011",
11921 => "010000110100001101000011",
11922 => "010000110100001101000011",
11923 => "010000110100001101000011",
11924 => "010000110100001101000011",
11925 => "010000110100001101000011",
11926 => "010000110100001101000011",
11927 => "010000110100001101000011",
11928 => "010000110100001101000011",
11929 => "010011100100111001001110",
11930 => "011001100110011001100110",
11931 => "011001100110011001100110",
11932 => "010000110100001101000011",
11933 => "010000110100001101000011",
11934 => "010000110100001101000011",
11935 => "010000110100001101000011",
11936 => "010000110100001101000011",
11937 => "010000110100001101000011",
11938 => "010000110100001101000011",
11939 => "010000110100001101000011",
11940 => "010000110100001101000011",
11941 => "001010000010100000101000",
11942 => "000101010001010100010101",
11943 => "000110000001100000011000",
11944 => "001000000010000000100000",
11945 => "001000000010000000100000",
11946 => "000000010000000100000001",
11947 => "000000000000000000000000",
11948 => "000000000000000000000000",
11949 => "000000000000000000000000",
11950 => "000000000000000000000000",
11951 => "000000000000000000000000",
11952 => "000000000000000000000000",
11953 => "000000000000000000000000",
11954 => "000000000000000000000000",
11955 => "000000000000000000000000",
11956 => "000000000000000000000000",
11957 => "000000000000000000000000",
11958 => "000000000000000000000000",
11959 => "000000000000000000000000",
11960 => "000000000000000000000000",
11961 => "000000000000000000000000",
11962 => "000000000000000000000000",
11963 => "000000000000000000000000",
11964 => "000000000000000000000000",
11965 => "000000000000000000000000",
11966 => "000000000000000000000000",
11967 => "000000000000000000000000",
11968 => "000000000000000000000000",
11969 => "000000000000000000000000",
11970 => "000000000000000000000000",
11971 => "000000000000000000000000",
11972 => "000000000000000000000000",
11973 => "000000000000000000000000",
11974 => "000000000000000000000000",
11975 => "000000000000000000000000",
11976 => "000000000000000000000000",
11977 => "000000000000000000000000",
11978 => "000000000000000000000000",
11979 => "000000000000000000000000",
11980 => "000000000000000000000000",
11981 => "000000000000000000000000",
11982 => "000000000000000000000000",
11983 => "000000000000000000000000",
11984 => "000000000000000000000000",
11985 => "000000000000000000000000",
11986 => "000000000000000000000000",
11987 => "000000000000000000000000",
11988 => "000000000000000000000000",
11989 => "000000000000000000000000",
11990 => "000000000000000000000000",
11991 => "000000000000000000000000",
11992 => "000000000000000000000000",
11993 => "000000000000000000000000",
11994 => "000000000000000000000000",
11995 => "000000000000000000000000",
11996 => "000000000000000000000000",
11997 => "000000000000000000000000",
11998 => "000000000000000000000000",
11999 => "000000000000000000000000",
12000 => "000000000000000000000000",
12001 => "000000000000000000000000",
12002 => "000000000000000000000000",
12003 => "000000000000000000000000",
12004 => "000000000000000000000000",
12005 => "000000000000000000000000",
12006 => "000000000000000000000000",
12007 => "000000000000000000000000",
12008 => "000000000000000000000000",
12009 => "000000000000000000000000",
12010 => "000000000000000000000000",
12011 => "000000000000000000000000",
12012 => "000000000000000000000000",
12013 => "000000000000000000000000",
12014 => "000000000000000000000000",
12015 => "000000000000000000000000",
12016 => "000000000000000000000000",
12017 => "000000000000000000000000",
12018 => "000000000000000000000000",
12019 => "000000000000000000000000",
12020 => "000000000000000000000000",
12021 => "000000000000000000000000",
12022 => "000000000000000000000000",
12023 => "000000000000000000000000",
12024 => "000000000000000000000000",
12025 => "000000000000000000000000",
12026 => "000000000000000000000000",
12027 => "000000000000000000000000",
12028 => "000000000000000000000000",
12029 => "000000000000000000000000",
12030 => "000000000000000000000000",
12031 => "000000000000000000000000",
12032 => "000000000000000000000000",
12033 => "000000000000000000000000",
12034 => "000000000000000000000000",
12035 => "000000000000000000000000",
12036 => "000000000000000000000000",
12037 => "000000000000000000000000",
12038 => "000000000000000000000000",
12039 => "000000000000000000000000",
12040 => "000000000000000000000000",
12041 => "000000000000000000000000",
12042 => "010110100101101001011010",
12043 => "011001100110011001100110",
12044 => "010101100101011001010110",
12045 => "010000110100001101000011",
12046 => "010000110100001101000011",
12047 => "010000110100001101000011",
12048 => "010000110100001101000011",
12049 => "010000110100001101000011",
12050 => "010000110100001101000011",
12051 => "010000110100001101000011",
12052 => "010000110100001101000011",
12053 => "010000110100001101000011",
12054 => "010000110100001101000011",
12055 => "010000110100001101000011",
12056 => "010111110101111101011111",
12057 => "011001100110011001100110",
12058 => "010110000101100001011000",
12059 => "010000110100001101000011",
12060 => "010000110100001101000011",
12061 => "010000110100001101000011",
12062 => "010000110100001101000011",
12063 => "010000110100001101000011",
12064 => "010000110100001101000011",
12065 => "010000110100001101000011",
12066 => "010000110100001101000011",
12067 => "010000110100001101000011",
12068 => "010000110100001101000011",
12069 => "010000110100001101000011",
12070 => "010000110100001101000011",
12071 => "010000110100001101000011",
12072 => "010000110100001101000011",
12073 => "010000110100001101000011",
12074 => "010000110100001101000011",
12075 => "010000110100001101000011",
12076 => "010000110100001101000011",
12077 => "010000110100001101000011",
12078 => "010000110100001101000011",
12079 => "010011100100111001001110",
12080 => "011001100110011001100110",
12081 => "011001100110011001100110",
12082 => "010000110100001101000011",
12083 => "010000110100001101000011",
12084 => "010000110100001101000011",
12085 => "010000110100001101000011",
12086 => "010000110100001101000011",
12087 => "010000110100001101000011",
12088 => "010000110100001101000011",
12089 => "010000110100001101000011",
12090 => "010000110100001101000011",
12091 => "010000110100001101000011",
12092 => "010000110100001101000011",
12093 => "010011000100110001001100",
12094 => "011001100110011001100110",
12095 => "011001100110011001100110",
12096 => "000000110000001100000011",
12097 => "000000000000000000000000",
12098 => "000000000000000000000000",
12099 => "000000000000000000000000",
12100 => "000000000000000000000000",
12101 => "000000000000000000000000",
12102 => "000000000000000000000000",
12103 => "000000000000000000000000",
12104 => "000000000000000000000000",
12105 => "000000000000000000000000",
12106 => "000000000000000000000000",
12107 => "000000000000000000000000",
12108 => "000000000000000000000000",
12109 => "000000000000000000000000",
12110 => "000000000000000000000000",
12111 => "000000000000000000000000",
12112 => "000000000000000000000000",
12113 => "000000000000000000000000",
12114 => "000000000000000000000000",
12115 => "000000000000000000000000",
12116 => "000000000000000000000000",
12117 => "000000000000000000000000",
12118 => "000000000000000000000000",
12119 => "000000000000000000000000",
12120 => "000000000000000000000000",
12121 => "000000000000000000000000",
12122 => "000000000000000000000000",
12123 => "000000000000000000000000",
12124 => "000000000000000000000000",
12125 => "000000000000000000000000",
12126 => "000000000000000000000000",
12127 => "000000000000000000000000",
12128 => "000000000000000000000000",
12129 => "000000000000000000000000",
12130 => "000000000000000000000000",
12131 => "000000000000000000000000",
12132 => "000000000000000000000000",
12133 => "000000000000000000000000",
12134 => "000000000000000000000000",
12135 => "000000000000000000000000",
12136 => "000000000000000000000000",
12137 => "000000000000000000000000",
12138 => "000000000000000000000000",
12139 => "000000000000000000000000",
12140 => "000000000000000000000000",
12141 => "000000000000000000000000",
12142 => "000000000000000000000000",
12143 => "000000000000000000000000",
12144 => "000000000000000000000000",
12145 => "000000000000000000000000",
12146 => "000000000000000000000000",
12147 => "000000000000000000000000",
12148 => "000000000000000000000000",
12149 => "000000000000000000000000",
12150 => "000000000000000000000000",
12151 => "000000000000000000000000",
12152 => "000000000000000000000000",
12153 => "000000000000000000000000",
12154 => "000000000000000000000000",
12155 => "000000000000000000000000",
12156 => "000000000000000000000000",
12157 => "000000000000000000000000",
12158 => "000000000000000000000000",
12159 => "000000000000000000000000",
12160 => "000000000000000000000000",
12161 => "000000000000000000000000",
12162 => "000000000000000000000000",
12163 => "000000000000000000000000",
12164 => "000000000000000000000000",
12165 => "000000000000000000000000",
12166 => "000000000000000000000000",
12167 => "000000000000000000000000",
12168 => "000000000000000000000000",
12169 => "000000000000000000000000",
12170 => "000000000000000000000000",
12171 => "000000000000000000000000",
12172 => "000000000000000000000000",
12173 => "000000000000000000000000",
12174 => "000000000000000000000000",
12175 => "000000000000000000000000",
12176 => "000000000000000000000000",
12177 => "000000000000000000000000",
12178 => "000000000000000000000000",
12179 => "000000000000000000000000",
12180 => "000000000000000000000000",
12181 => "000000000000000000000000",
12182 => "000000000000000000000000",
12183 => "000000000000000000000000",
12184 => "000000000000000000000000",
12185 => "000000000000000000000000",
12186 => "000000000000000000000000",
12187 => "000000000000000000000000",
12188 => "000000000000000000000000",
12189 => "000000000000000000000000",
12190 => "000000000000000000000000",
12191 => "000000000000000000000000",
12192 => "010110100101101001011010",
12193 => "011001100110011001100110",
12194 => "010101100101011001010110",
12195 => "010000110100001101000011",
12196 => "010000110100001101000011",
12197 => "010000110100001101000011",
12198 => "010000110100001101000011",
12199 => "010000110100001101000011",
12200 => "010000110100001101000011",
12201 => "010000110100001101000011",
12202 => "010000110100001101000011",
12203 => "010000110100001101000011",
12204 => "010000110100001101000011",
12205 => "010000110100001101000011",
12206 => "010111110101111101011111",
12207 => "011001100110011001100110",
12208 => "010110000101100001011000",
12209 => "010000110100001101000011",
12210 => "010000110100001101000011",
12211 => "010000110100001101000011",
12212 => "010000110100001101000011",
12213 => "010000110100001101000011",
12214 => "010000110100001101000011",
12215 => "010000110100001101000011",
12216 => "010000110100001101000011",
12217 => "010000110100001101000011",
12218 => "010000110100001101000011",
12219 => "010000110100001101000011",
12220 => "010000110100001101000011",
12221 => "010000110100001101000011",
12222 => "010000110100001101000011",
12223 => "010000110100001101000011",
12224 => "010000110100001101000011",
12225 => "010000110100001101000011",
12226 => "010000110100001101000011",
12227 => "010000110100001101000011",
12228 => "010000110100001101000011",
12229 => "010011100100111001001110",
12230 => "011001100110011001100110",
12231 => "011001100110011001100110",
12232 => "010000110100001101000011",
12233 => "010000110100001101000011",
12234 => "010000110100001101000011",
12235 => "010000110100001101000011",
12236 => "010000110100001101000011",
12237 => "010000110100001101000011",
12238 => "010000110100001101000011",
12239 => "010000110100001101000011",
12240 => "010000110100001101000011",
12241 => "010000110100001101000011",
12242 => "010000110100001101000011",
12243 => "010011000100110001001100",
12244 => "011001100110011001100110",
12245 => "011001100110011001100110",
12246 => "000000110000001100000011",
12247 => "000000000000000000000000",
12248 => "000000000000000000000000",
12249 => "000000000000000000000000",
12250 => "000000000000000000000000",
12251 => "000000000000000000000000",
12252 => "000000000000000000000000",
12253 => "000000000000000000000000",
12254 => "000000000000000000000000",
12255 => "000000000000000000000000",
12256 => "000000000000000000000000",
12257 => "000000000000000000000000",
12258 => "000000000000000000000000",
12259 => "000000000000000000000000",
12260 => "000000000000000000000000",
12261 => "000000000000000000000000",
12262 => "000000000000000000000000",
12263 => "000000000000000000000000",
12264 => "000000000000000000000000",
12265 => "000000000000000000000000",
12266 => "000000000000000000000000",
12267 => "000000000000000000000000",
12268 => "000000000000000000000000",
12269 => "000000000000000000000000",
12270 => "000000000000000000000000",
12271 => "000000000000000000000000",
12272 => "000000000000000000000000",
12273 => "000000000000000000000000",
12274 => "000000000000000000000000",
12275 => "000000000000000000000000",
12276 => "000000000000000000000000",
12277 => "000000000000000000000000",
12278 => "000000000000000000000000",
12279 => "000000000000000000000000",
12280 => "000000000000000000000000",
12281 => "000000000000000000000000",
12282 => "000000000000000000000000",
12283 => "000000000000000000000000",
12284 => "000000000000000000000000",
12285 => "000000000000000000000000",
12286 => "000000000000000000000000",
12287 => "000000000000000000000000",
12288 => "000000000000000000000000",
12289 => "000000000000000000000000",
12290 => "000000000000000000000000",
12291 => "000000000000000000000000",
12292 => "000000000000000000000000",
12293 => "000000000000000000000000",
12294 => "000000000000000000000000",
12295 => "000000000000000000000000",
12296 => "000000000000000000000000",
12297 => "000000000000000000000000",
12298 => "000000000000000000000000",
12299 => "000000000000000000000000",
12300 => "000000000000000000000000",
12301 => "000000000000000000000000",
12302 => "000000000000000000000000",
12303 => "000000000000000000000000",
12304 => "000000000000000000000000",
12305 => "000000000000000000000000",
12306 => "000000000000000000000000",
12307 => "000000000000000000000000",
12308 => "000000000000000000000000",
12309 => "000000000000000000000000",
12310 => "000000000000000000000000",
12311 => "000000000000000000000000",
12312 => "000000000000000000000000",
12313 => "000000000000000000000000",
12314 => "000000000000000000000000",
12315 => "000000000000000000000000",
12316 => "000000000000000000000000",
12317 => "000000000000000000000000",
12318 => "000000000000000000000000",
12319 => "000000000000000000000000",
12320 => "000000000000000000000000",
12321 => "000000000000000000000000",
12322 => "000000000000000000000000",
12323 => "000000000000000000000000",
12324 => "000000000000000000000000",
12325 => "000000000000000000000000",
12326 => "000000000000000000000000",
12327 => "000000000000000000000000",
12328 => "000000000000000000000000",
12329 => "000000000000000000000000",
12330 => "000000000000000000000000",
12331 => "000000000000000000000000",
12332 => "000000000000000000000000",
12333 => "000000000000000000000000",
12334 => "000000000000000000000000",
12335 => "000000000000000000000000",
12336 => "000000000000000000000000",
12337 => "000000000000000000000000",
12338 => "000000000000000000000000",
12339 => "000010100000101000001010",
12340 => "010000110100001101000011",
12341 => "010000110100001101000011",
12342 => "011000100110001001100010",
12343 => "011001100110011001100110",
12344 => "010101100101011001010110",
12345 => "010000110100001101000011",
12346 => "010000110100001101000011",
12347 => "010000110100001101000011",
12348 => "010000110100001101000011",
12349 => "010000110100001101000011",
12350 => "010000110100001101000011",
12351 => "010000110100001101000011",
12352 => "010000110100001101000011",
12353 => "010000110100001101000011",
12354 => "010000110100001101000011",
12355 => "010000110100001101000011",
12356 => "010111110101111101011111",
12357 => "011001100110011001100110",
12358 => "010110000101100001011000",
12359 => "010000110100001101000011",
12360 => "010000110100001101000011",
12361 => "010000110100001101000011",
12362 => "010000110100001101000011",
12363 => "010000110100001101000011",
12364 => "010000110100001101000011",
12365 => "010000110100001101000011",
12366 => "010000110100001101000011",
12367 => "010000110100001101000011",
12368 => "010000110100001101000011",
12369 => "010000110100001101000011",
12370 => "010000110100001101000011",
12371 => "010000110100001101000011",
12372 => "010000110100001101000011",
12373 => "010000110100001101000011",
12374 => "010000110100001101000011",
12375 => "010000110100001101000011",
12376 => "010000110100001101000011",
12377 => "010000110100001101000011",
12378 => "010000110100001101000011",
12379 => "010011100100111001001110",
12380 => "011001100110011001100110",
12381 => "011001100110011001100110",
12382 => "010000110100001101000011",
12383 => "010000110100001101000011",
12384 => "010000110100001101000011",
12385 => "010000110100001101000011",
12386 => "010000110100001101000011",
12387 => "010000110100001101000011",
12388 => "010000110100001101000011",
12389 => "010000110100001101000011",
12390 => "010000110100001101000011",
12391 => "010000110100001101000011",
12392 => "010000110100001101000011",
12393 => "010011000100110001001100",
12394 => "011001100110011001100110",
12395 => "011001100110011001100110",
12396 => "010001000100010001000100",
12397 => "010000110100001101000011",
12398 => "000111010001110100011101",
12399 => "000000000000000000000000",
12400 => "000000000000000000000000",
12401 => "000000000000000000000000",
12402 => "000000000000000000000000",
12403 => "000000000000000000000000",
12404 => "000000000000000000000000",
12405 => "000000000000000000000000",
12406 => "000000000000000000000000",
12407 => "000000000000000000000000",
12408 => "000000000000000000000000",
12409 => "000000000000000000000000",
12410 => "000000000000000000000000",
12411 => "000000000000000000000000",
12412 => "000000000000000000000000",
12413 => "000000000000000000000000",
12414 => "000000000000000000000000",
12415 => "000000000000000000000000",
12416 => "000000000000000000000000",
12417 => "000000000000000000000000",
12418 => "000000000000000000000000",
12419 => "000000000000000000000000",
12420 => "000000000000000000000000",
12421 => "000000000000000000000000",
12422 => "000000000000000000000000",
12423 => "000000000000000000000000",
12424 => "000000000000000000000000",
12425 => "000000000000000000000000",
12426 => "000000000000000000000000",
12427 => "000000000000000000000000",
12428 => "000000000000000000000000",
12429 => "000000000000000000000000",
12430 => "000000000000000000000000",
12431 => "000000000000000000000000",
12432 => "000000000000000000000000",
12433 => "000000000000000000000000",
12434 => "000000000000000000000000",
12435 => "000000000000000000000000",
12436 => "000000000000000000000000",
12437 => "000000000000000000000000",
12438 => "000000000000000000000000",
12439 => "000000000000000000000000",
12440 => "000000000000000000000000",
12441 => "000000000000000000000000",
12442 => "000000000000000000000000",
12443 => "000000000000000000000000",
12444 => "000000000000000000000000",
12445 => "000000000000000000000000",
12446 => "000000000000000000000000",
12447 => "000000000000000000000000",
12448 => "000000000000000000000000",
12449 => "000000000000000000000000",
12450 => "000000000000000000000000",
12451 => "000000000000000000000000",
12452 => "000000000000000000000000",
12453 => "000000000000000000000000",
12454 => "000000000000000000000000",
12455 => "000000000000000000000000",
12456 => "000000000000000000000000",
12457 => "000000000000000000000000",
12458 => "000000000000000000000000",
12459 => "000000000000000000000000",
12460 => "000000000000000000000000",
12461 => "000000000000000000000000",
12462 => "000000000000000000000000",
12463 => "000000000000000000000000",
12464 => "000000000000000000000000",
12465 => "000000000000000000000000",
12466 => "000000000000000000000000",
12467 => "000000000000000000000000",
12468 => "000000000000000000000000",
12469 => "000000000000000000000000",
12470 => "000000000000000000000000",
12471 => "000000000000000000000000",
12472 => "000000000000000000000000",
12473 => "000000000000000000000000",
12474 => "000000000000000000000000",
12475 => "000000000000000000000000",
12476 => "000000000000000000000000",
12477 => "000000000000000000000000",
12478 => "000000000000000000000000",
12479 => "000000000000000000000000",
12480 => "000000000000000000000000",
12481 => "000000000000000000000000",
12482 => "000000000000000000000000",
12483 => "000000000000000000000000",
12484 => "000000000000000000000000",
12485 => "000000000000000000000000",
12486 => "000000000000000000000000",
12487 => "000000000000000000000000",
12488 => "000000000000000000000000",
12489 => "000010100000101000001010",
12490 => "010000110100001101000011",
12491 => "010000110100001101000011",
12492 => "011000100110001001100010",
12493 => "011001100110011001100110",
12494 => "010101100101011001010110",
12495 => "010000110100001101000011",
12496 => "010000110100001101000011",
12497 => "010000110100001101000011",
12498 => "010000110100001101000011",
12499 => "010000110100001101000011",
12500 => "010000110100001101000011",
12501 => "010000110100001101000011",
12502 => "010000110100001101000011",
12503 => "010000110100001101000011",
12504 => "010000110100001101000011",
12505 => "010000110100001101000011",
12506 => "010111110101111101011111",
12507 => "011001100110011001100110",
12508 => "010110000101100001011000",
12509 => "010000110100001101000011",
12510 => "010000110100001101000011",
12511 => "010000110100001101000011",
12512 => "010000110100001101000011",
12513 => "010000110100001101000011",
12514 => "010000110100001101000011",
12515 => "010000110100001101000011",
12516 => "010000110100001101000011",
12517 => "010000110100001101000011",
12518 => "010000110100001101000011",
12519 => "010000110100001101000011",
12520 => "010000110100001101000011",
12521 => "010000110100001101000011",
12522 => "010000110100001101000011",
12523 => "010000110100001101000011",
12524 => "010000110100001101000011",
12525 => "010000110100001101000011",
12526 => "010000110100001101000011",
12527 => "010000110100001101000011",
12528 => "010000110100001101000011",
12529 => "010011100100111001001110",
12530 => "011001100110011001100110",
12531 => "011001100110011001100110",
12532 => "010000110100001101000011",
12533 => "010000110100001101000011",
12534 => "010000110100001101000011",
12535 => "010000110100001101000011",
12536 => "010000110100001101000011",
12537 => "010000110100001101000011",
12538 => "010000110100001101000011",
12539 => "010000110100001101000011",
12540 => "010000110100001101000011",
12541 => "010000110100001101000011",
12542 => "010000110100001101000011",
12543 => "010011000100110001001100",
12544 => "011001100110011001100110",
12545 => "011001100110011001100110",
12546 => "010001000100010001000100",
12547 => "010000110100001101000011",
12548 => "000111010001110100011101",
12549 => "000000000000000000000000",
12550 => "000000000000000000000000",
12551 => "000000000000000000000000",
12552 => "000000000000000000000000",
12553 => "000000000000000000000000",
12554 => "000000000000000000000000",
12555 => "000000000000000000000000",
12556 => "000000000000000000000000",
12557 => "000000000000000000000000",
12558 => "000000000000000000000000",
12559 => "000000000000000000000000",
12560 => "000000000000000000000000",
12561 => "000000000000000000000000",
12562 => "000000000000000000000000",
12563 => "000000000000000000000000",
12564 => "000000000000000000000000",
12565 => "000000000000000000000000",
12566 => "000000000000000000000000",
12567 => "000000000000000000000000",
12568 => "000000000000000000000000",
12569 => "000000000000000000000000",
12570 => "000000000000000000000000",
12571 => "000000000000000000000000",
12572 => "000000000000000000000000",
12573 => "000000000000000000000000",
12574 => "000000000000000000000000",
12575 => "000000000000000000000000",
12576 => "000000000000000000000000",
12577 => "000000000000000000000000",
12578 => "000000000000000000000000",
12579 => "000000000000000000000000",
12580 => "000000000000000000000000",
12581 => "000000000000000000000000",
12582 => "000000000000000000000000",
12583 => "000000000000000000000000",
12584 => "000000000000000000000000",
12585 => "000000000000000000000000",
12586 => "000000000000000000000000",
12587 => "000000000000000000000000",
12588 => "000000000000000000000000",
12589 => "000000000000000000000000",
12590 => "000000000000000000000000",
12591 => "000000000000000000000000",
12592 => "000000000000000000000000",
12593 => "000000000000000000000000",
12594 => "000000000000000000000000",
12595 => "000000000000000000000000",
12596 => "000000000000000000000000",
12597 => "000000000000000000000000",
12598 => "000000000000000000000000",
12599 => "000000000000000000000000",
12600 => "000000000000000000000000",
12601 => "000000000000000000000000",
12602 => "000000000000000000000000",
12603 => "000000000000000000000000",
12604 => "000000000000000000000000",
12605 => "000000000000000000000000",
12606 => "000000000000000000000000",
12607 => "000000000000000000000000",
12608 => "000000000000000000000000",
12609 => "000000000000000000000000",
12610 => "000000000000000000000000",
12611 => "000000000000000000000000",
12612 => "000000000000000000000000",
12613 => "000000000000000000000000",
12614 => "000000000000000000000000",
12615 => "000000000000000000000000",
12616 => "000000000000000000000000",
12617 => "000000000000000000000000",
12618 => "000000000000000000000000",
12619 => "000000000000000000000000",
12620 => "000000000000000000000000",
12621 => "000000000000000000000000",
12622 => "000000000000000000000000",
12623 => "000000000000000000000000",
12624 => "000000000000000000000000",
12625 => "000000000000000000000000",
12626 => "000000000000000000000000",
12627 => "000000000000000000000000",
12628 => "000000000000000000000000",
12629 => "000000000000000000000000",
12630 => "000000000000000000000000",
12631 => "000000000000000000000000",
12632 => "000000000000000000000000",
12633 => "000000000000000000000000",
12634 => "000000000000000000000000",
12635 => "001001100010011000100110",
12636 => "001010100010101000101010",
12637 => "001010100010101000101010",
12638 => "001010100010101000101010",
12639 => "001100010011000100110001",
12640 => "010110010101100101011001",
12641 => "010110010101100101011001",
12642 => "010100010101000101010001",
12643 => "010100000101000001010000",
12644 => "010010100100101001001010",
12645 => "010000110100001101000011",
12646 => "010001100100011001000110",
12647 => "010110010101100101011001",
12648 => "010110010101100101011001",
12649 => "010001110100011101000111",
12650 => "010000110100001101000011",
12651 => "010000110100001101000011",
12652 => "010000110100001101000011",
12653 => "010000110100001101000011",
12654 => "010000110100001101000011",
12655 => "010000110100001101000011",
12656 => "010011010100110101001101",
12657 => "010100000101000001010000",
12658 => "010010110100101101001011",
12659 => "010000110100001101000011",
12660 => "010000110100001101000011",
12661 => "010000110100001101000011",
12662 => "010000110100001101000011",
12663 => "010000110100001101000011",
12664 => "010000110100001101000011",
12665 => "010000110100001101000011",
12666 => "010000110100001101000011",
12667 => "010000110100001101000011",
12668 => "010000110100001101000011",
12669 => "010000110100001101000011",
12670 => "010000110100001101000011",
12671 => "010000110100001101000011",
12672 => "010000110100001101000011",
12673 => "010000110100001101000011",
12674 => "010000110100001101000011",
12675 => "010000110100001101000011",
12676 => "010000110100001101000011",
12677 => "010000110100001101000011",
12678 => "010000110100001101000011",
12679 => "010001110100011101000111",
12680 => "010100000101000001010000",
12681 => "010100000101000001010000",
12682 => "010000110100001101000011",
12683 => "010000110100001101000011",
12684 => "010000110100001101000011",
12685 => "010000110100001101000011",
12686 => "010000110100001101000011",
12687 => "010000110100001101000011",
12688 => "010000110100001101000011",
12689 => "010110010101100101011001",
12690 => "010110010101100101011001",
12691 => "010011000100110001001100",
12692 => "010000110100001101000011",
12693 => "010001100100011001000110",
12694 => "010100000101000001010000",
12695 => "010100000101000001010000",
12696 => "010110010101100101011001",
12697 => "010110010101100101011001",
12698 => "001111100011111000111110",
12699 => "001010100010101000101010",
12700 => "001010100010101000101010",
12701 => "001010100010101000101010",
12702 => "001010100010101000101010",
12703 => "000000100000001000000010",
12704 => "000000000000000000000000",
12705 => "000000000000000000000000",
12706 => "000000000000000000000000",
12707 => "000000000000000000000000",
12708 => "000000000000000000000000",
12709 => "000000000000000000000000",
12710 => "000000000000000000000000",
12711 => "000000000000000000000000",
12712 => "000000000000000000000000",
12713 => "000000000000000000000000",
12714 => "000000000000000000000000",
12715 => "000000000000000000000000",
12716 => "000000000000000000000000",
12717 => "000000000000000000000000",
12718 => "000000000000000000000000",
12719 => "000000000000000000000000",
12720 => "000000000000000000000000",
12721 => "000000000000000000000000",
12722 => "000000000000000000000000",
12723 => "000000000000000000000000",
12724 => "000000000000000000000000",
12725 => "000000000000000000000000",
12726 => "000000000000000000000000",
12727 => "000000000000000000000000",
12728 => "000000000000000000000000",
12729 => "000000000000000000000000",
12730 => "000000000000000000000000",
12731 => "000000000000000000000000",
12732 => "000000000000000000000000",
12733 => "000000000000000000000000",
12734 => "000000000000000000000000",
12735 => "000000000000000000000000",
12736 => "000000000000000000000000",
12737 => "000000000000000000000000",
12738 => "000000000000000000000000",
12739 => "000000000000000000000000",
12740 => "000000000000000000000000",
12741 => "000000000000000000000000",
12742 => "000000000000000000000000",
12743 => "000000000000000000000000",
12744 => "000000000000000000000000",
12745 => "000000000000000000000000",
12746 => "000000000000000000000000",
12747 => "000000000000000000000000",
12748 => "000000000000000000000000",
12749 => "000000000000000000000000",
12750 => "000000000000000000000000",
12751 => "000000000000000000000000",
12752 => "000000000000000000000000",
12753 => "000000000000000000000000",
12754 => "000000000000000000000000",
12755 => "000000000000000000000000",
12756 => "000000000000000000000000",
12757 => "000000000000000000000000",
12758 => "000000000000000000000000",
12759 => "000000000000000000000000",
12760 => "000000000000000000000000",
12761 => "000000000000000000000000",
12762 => "000000000000000000000000",
12763 => "000000000000000000000000",
12764 => "000000000000000000000000",
12765 => "000000000000000000000000",
12766 => "000000000000000000000000",
12767 => "000000000000000000000000",
12768 => "000000000000000000000000",
12769 => "000000000000000000000000",
12770 => "000000000000000000000000",
12771 => "000000000000000000000000",
12772 => "000000000000000000000000",
12773 => "000000000000000000000000",
12774 => "000000000000000000000000",
12775 => "000000000000000000000000",
12776 => "000000000000000000000000",
12777 => "000000000000000000000000",
12778 => "000000000000000000000000",
12779 => "000000000000000000000000",
12780 => "000000000000000000000000",
12781 => "000000000000000000000000",
12782 => "000000000000000000000000",
12783 => "000000000000000000000000",
12784 => "000000000000000000000000",
12785 => "001111010011110100111101",
12786 => "010000110100001101000011",
12787 => "010000110100001101000011",
12788 => "010000110100001101000011",
12789 => "010010000100100001001000",
12790 => "011001100110011001100110",
12791 => "011001100110011001100110",
12792 => "010001110100011101000111",
12793 => "010000110100001101000011",
12794 => "010000110100001101000011",
12795 => "010000110100001101000011",
12796 => "010001110100011101000111",
12797 => "011001100110011001100110",
12798 => "011001100110011001100110",
12799 => "010010010100100101001001",
12800 => "010000110100001101000011",
12801 => "010000110100001101000011",
12802 => "010000110100001101000011",
12803 => "010000110100001101000011",
12804 => "010000110100001101000011",
12805 => "010000110100001101000011",
12806 => "010000110100001101000011",
12807 => "010000110100001101000011",
12808 => "010000110100001101000011",
12809 => "010000110100001101000011",
12810 => "010000110100001101000011",
12811 => "010000110100001101000011",
12812 => "010000110100001101000011",
12813 => "010000110100001101000011",
12814 => "010000110100001101000011",
12815 => "010000110100001101000011",
12816 => "010000110100001101000011",
12817 => "010000110100001101000011",
12818 => "010000110100001101000011",
12819 => "010000110100001101000011",
12820 => "010000110100001101000011",
12821 => "010000110100001101000011",
12822 => "010000110100001101000011",
12823 => "010000110100001101000011",
12824 => "010000110100001101000011",
12825 => "010000110100001101000011",
12826 => "010000110100001101000011",
12827 => "010000110100001101000011",
12828 => "010000110100001101000011",
12829 => "010000110100001101000011",
12830 => "010000110100001101000011",
12831 => "010000110100001101000011",
12832 => "010000110100001101000011",
12833 => "010000110100001101000011",
12834 => "010000110100001101000011",
12835 => "010000110100001101000011",
12836 => "010000110100001101000011",
12837 => "010000110100001101000011",
12838 => "010000110100001101000011",
12839 => "011001100110011001100110",
12840 => "011001100110011001100110",
12841 => "010100010101000101010001",
12842 => "010000110100001101000011",
12843 => "010000110100001101000011",
12844 => "010000110100001101000011",
12845 => "010000110100001101000011",
12846 => "011001010110010101100101",
12847 => "011001100110011001100110",
12848 => "010100100101001001010010",
12849 => "010000110100001101000011",
12850 => "010000110100001101000011",
12851 => "010000110100001101000011",
12852 => "010000110100001101000011",
12853 => "000001000000010000000100",
12854 => "000000000000000000000000",
12855 => "000000000000000000000000",
12856 => "000000000000000000000000",
12857 => "000000000000000000000000",
12858 => "000000000000000000000000",
12859 => "000000000000000000000000",
12860 => "000000000000000000000000",
12861 => "000000000000000000000000",
12862 => "000000000000000000000000",
12863 => "000000000000000000000000",
12864 => "000000000000000000000000",
12865 => "000000000000000000000000",
12866 => "000000000000000000000000",
12867 => "000000000000000000000000",
12868 => "000000000000000000000000",
12869 => "000000000000000000000000",
12870 => "000000000000000000000000",
12871 => "000000000000000000000000",
12872 => "000000000000000000000000",
12873 => "000000000000000000000000",
12874 => "000000000000000000000000",
12875 => "000000000000000000000000",
12876 => "000000000000000000000000",
12877 => "000000000000000000000000",
12878 => "000000000000000000000000",
12879 => "000000000000000000000000",
12880 => "000000000000000000000000",
12881 => "000000000000000000000000",
12882 => "000000000000000000000000",
12883 => "000000000000000000000000",
12884 => "000000000000000000000000",
12885 => "000000000000000000000000",
12886 => "000000000000000000000000",
12887 => "000000000000000000000000",
12888 => "000000000000000000000000",
12889 => "000000000000000000000000",
12890 => "000000000000000000000000",
12891 => "000000000000000000000000",
12892 => "000000000000000000000000",
12893 => "000000000000000000000000",
12894 => "000000000000000000000000",
12895 => "000000000000000000000000",
12896 => "000000000000000000000000",
12897 => "000000000000000000000000",
12898 => "000000000000000000000000",
12899 => "000000000000000000000000",
12900 => "000000000000000000000000",
12901 => "000000000000000000000000",
12902 => "000000000000000000000000",
12903 => "000000000000000000000000",
12904 => "000000000000000000000000",
12905 => "000000000000000000000000",
12906 => "000000000000000000000000",
12907 => "000000000000000000000000",
12908 => "000000000000000000000000",
12909 => "000000000000000000000000",
12910 => "000000000000000000000000",
12911 => "000000000000000000000000",
12912 => "000000000000000000000000",
12913 => "000000000000000000000000",
12914 => "000000000000000000000000",
12915 => "000000000000000000000000",
12916 => "000000000000000000000000",
12917 => "000000000000000000000000",
12918 => "000000000000000000000000",
12919 => "000000000000000000000000",
12920 => "000000000000000000000000",
12921 => "000000000000000000000000",
12922 => "000000000000000000000000",
12923 => "000000000000000000000000",
12924 => "000000000000000000000000",
12925 => "000000000000000000000000",
12926 => "000000000000000000000000",
12927 => "000000000000000000000000",
12928 => "000000000000000000000000",
12929 => "000000000000000000000000",
12930 => "000000000000000000000000",
12931 => "000000000000000000000000",
12932 => "000001000000010000000100",
12933 => "000100110001001100010011",
12934 => "000100110001001100010011",
12935 => "010010000100100001001000",
12936 => "010011010100110101001101",
12937 => "010011010100110101001101",
12938 => "010011010100110101001101",
12939 => "010011110100111101001111",
12940 => "010111000101110001011100",
12941 => "010111000101110001011100",
12942 => "010001100100011001000110",
12943 => "010000110100001101000011",
12944 => "010000110100001101000011",
12945 => "010000110100001101000011",
12946 => "010001110100011101000111",
12947 => "011001100110011001100110",
12948 => "011001100110011001100110",
12949 => "010010010100100101001001",
12950 => "010000110100001101000011",
12951 => "010000110100001101000011",
12952 => "010000110100001101000011",
12953 => "010000110100001101000011",
12954 => "010000110100001101000011",
12955 => "010000110100001101000011",
12956 => "010000110100001101000011",
12957 => "010000110100001101000011",
12958 => "010000110100001101000011",
12959 => "010000110100001101000011",
12960 => "010000110100001101000011",
12961 => "010000110100001101000011",
12962 => "010000110100001101000011",
12963 => "010000110100001101000011",
12964 => "010000110100001101000011",
12965 => "010000110100001101000011",
12966 => "010000110100001101000011",
12967 => "010000110100001101000011",
12968 => "010000110100001101000011",
12969 => "010000110100001101000011",
12970 => "010000110100001101000011",
12971 => "010000110100001101000011",
12972 => "010000110100001101000011",
12973 => "010000110100001101000011",
12974 => "010000110100001101000011",
12975 => "010000110100001101000011",
12976 => "010000110100001101000011",
12977 => "010000110100001101000011",
12978 => "010000110100001101000011",
12979 => "010000110100001101000011",
12980 => "010000110100001101000011",
12981 => "010000110100001101000011",
12982 => "010000110100001101000011",
12983 => "010000110100001101000011",
12984 => "010000110100001101000011",
12985 => "010000110100001101000011",
12986 => "010000110100001101000011",
12987 => "010000110100001101000011",
12988 => "010000110100001101000011",
12989 => "011001100110011001100110",
12990 => "011001100110011001100110",
12991 => "010100010101000101010001",
12992 => "010000110100001101000011",
12993 => "010000110100001101000011",
12994 => "010000110100001101000011",
12995 => "010000110100001101000011",
12996 => "010110110101101101011011",
12997 => "010111000101110001011100",
12998 => "010101000101010001010100",
12999 => "010011010100110101001101",
13000 => "010011010100110101001101",
13001 => "010011010100110101001101",
13002 => "010011010100110101001101",
13003 => "000101100001011000010110",
13004 => "000100110001001100010011",
13005 => "000010010000100100001001",
13006 => "000000000000000000000000",
13007 => "000000000000000000000000",
13008 => "000000000000000000000000",
13009 => "000000000000000000000000",
13010 => "000000000000000000000000",
13011 => "000000000000000000000000",
13012 => "000000000000000000000000",
13013 => "000000000000000000000000",
13014 => "000000000000000000000000",
13015 => "000000000000000000000000",
13016 => "000000000000000000000000",
13017 => "000000000000000000000000",
13018 => "000000000000000000000000",
13019 => "000000000000000000000000",
13020 => "000000000000000000000000",
13021 => "000000000000000000000000",
13022 => "000000000000000000000000",
13023 => "000000000000000000000000",
13024 => "000000000000000000000000",
13025 => "000000000000000000000000",
13026 => "000000000000000000000000",
13027 => "000000000000000000000000",
13028 => "000000000000000000000000",
13029 => "000000000000000000000000",
13030 => "000000000000000000000000",
13031 => "000000000000000000000000",
13032 => "000000000000000000000000",
13033 => "000000000000000000000000",
13034 => "000000000000000000000000",
13035 => "000000000000000000000000",
13036 => "000000000000000000000000",
13037 => "000000000000000000000000",
13038 => "000000000000000000000000",
13039 => "000000000000000000000000",
13040 => "000000000000000000000000",
13041 => "000000000000000000000000",
13042 => "000000000000000000000000",
13043 => "000000000000000000000000",
13044 => "000000000000000000000000",
13045 => "000000000000000000000000",
13046 => "000000000000000000000000",
13047 => "000000000000000000000000",
13048 => "000000000000000000000000",
13049 => "000000000000000000000000",
13050 => "000000000000000000000000",
13051 => "000000000000000000000000",
13052 => "000000000000000000000000",
13053 => "000000000000000000000000",
13054 => "000000000000000000000000",
13055 => "000000000000000000000000",
13056 => "000000000000000000000000",
13057 => "000000000000000000000000",
13058 => "000000000000000000000000",
13059 => "000000000000000000000000",
13060 => "000000000000000000000000",
13061 => "000000000000000000000000",
13062 => "000000000000000000000000",
13063 => "000000000000000000000000",
13064 => "000000000000000000000000",
13065 => "000000000000000000000000",
13066 => "000000000000000000000000",
13067 => "000000000000000000000000",
13068 => "000000000000000000000000",
13069 => "000000000000000000000000",
13070 => "000000000000000000000000",
13071 => "000000000000000000000000",
13072 => "000000000000000000000000",
13073 => "000000000000000000000000",
13074 => "000000000000000000000000",
13075 => "000000000000000000000000",
13076 => "000000000000000000000000",
13077 => "000000000000000000000000",
13078 => "000000000000000000000000",
13079 => "000000000000000000000000",
13080 => "000000000000000000000000",
13081 => "000000000000000000000000",
13082 => "000011010000110100001101",
13083 => "010000110100001101000011",
13084 => "010000110100001101000011",
13085 => "011000110110001101100011",
13086 => "011001100110011001100110",
13087 => "011001100110011001100110",
13088 => "011001100110011001100110",
13089 => "011000010110000101100001",
13090 => "010000110100001101000011",
13091 => "010000110100001101000011",
13092 => "010000110100001101000011",
13093 => "010000110100001101000011",
13094 => "010000110100001101000011",
13095 => "010000110100001101000011",
13096 => "010001110100011101000111",
13097 => "011001100110011001100110",
13098 => "011001100110011001100110",
13099 => "010010010100100101001001",
13100 => "010000110100001101000011",
13101 => "010000110100001101000011",
13102 => "010000110100001101000011",
13103 => "010000110100001101000011",
13104 => "010000110100001101000011",
13105 => "010000110100001101000011",
13106 => "010000110100001101000011",
13107 => "010000110100001101000011",
13108 => "010000110100001101000011",
13109 => "010000110100001101000011",
13110 => "010000110100001101000011",
13111 => "010000110100001101000011",
13112 => "010000110100001101000011",
13113 => "010000110100001101000011",
13114 => "010000110100001101000011",
13115 => "010000110100001101000011",
13116 => "010000110100001101000011",
13117 => "010000110100001101000011",
13118 => "010000110100001101000011",
13119 => "010000110100001101000011",
13120 => "010000110100001101000011",
13121 => "010000110100001101000011",
13122 => "010000110100001101000011",
13123 => "010000110100001101000011",
13124 => "010000110100001101000011",
13125 => "010000110100001101000011",
13126 => "010000110100001101000011",
13127 => "010000110100001101000011",
13128 => "010000110100001101000011",
13129 => "010000110100001101000011",
13130 => "010000110100001101000011",
13131 => "010000110100001101000011",
13132 => "010000110100001101000011",
13133 => "010000110100001101000011",
13134 => "010000110100001101000011",
13135 => "010000110100001101000011",
13136 => "010000110100001101000011",
13137 => "010000110100001101000011",
13138 => "010000110100001101000011",
13139 => "011001100110011001100110",
13140 => "011001100110011001100110",
13141 => "010100010101000101010001",
13142 => "010000110100001101000011",
13143 => "010000110100001101000011",
13144 => "010000110100001101000011",
13145 => "010000110100001101000011",
13146 => "010000110100001101000011",
13147 => "010000110100001101000011",
13148 => "010101110101011101010111",
13149 => "011001100110011001100110",
13150 => "011001100110011001100110",
13151 => "011001100110011001100110",
13152 => "011001100110011001100110",
13153 => "010001010100010101000101",
13154 => "010000110100001101000011",
13155 => "000111110001111100011111",
13156 => "000000000000000000000000",
13157 => "000000000000000000000000",
13158 => "000000000000000000000000",
13159 => "000000000000000000000000",
13160 => "000000000000000000000000",
13161 => "000000000000000000000000",
13162 => "000000000000000000000000",
13163 => "000000000000000000000000",
13164 => "000000000000000000000000",
13165 => "000000000000000000000000",
13166 => "000000000000000000000000",
13167 => "000000000000000000000000",
13168 => "000000000000000000000000",
13169 => "000000000000000000000000",
13170 => "000000000000000000000000",
13171 => "000000000000000000000000",
13172 => "000000000000000000000000",
13173 => "000000000000000000000000",
13174 => "000000000000000000000000",
13175 => "000000000000000000000000",
13176 => "000000000000000000000000",
13177 => "000000000000000000000000",
13178 => "000000000000000000000000",
13179 => "000000000000000000000000",
13180 => "000000000000000000000000",
13181 => "000000000000000000000000",
13182 => "000000000000000000000000",
13183 => "000000000000000000000000",
13184 => "000000000000000000000000",
13185 => "000000000000000000000000",
13186 => "000000000000000000000000",
13187 => "000000000000000000000000",
13188 => "000000000000000000000000",
13189 => "000000000000000000000000",
13190 => "000000000000000000000000",
13191 => "000000000000000000000000",
13192 => "000000000000000000000000",
13193 => "000000000000000000000000",
13194 => "000000000000000000000000",
13195 => "000000000000000000000000",
13196 => "000000000000000000000000",
13197 => "000000000000000000000000",
13198 => "000000000000000000000000",
13199 => "000000000000000000000000",
13200 => "000000000000000000000000",
13201 => "000000000000000000000000",
13202 => "000000000000000000000000",
13203 => "000000000000000000000000",
13204 => "000000000000000000000000",
13205 => "000000000000000000000000",
13206 => "000000000000000000000000",
13207 => "000000000000000000000000",
13208 => "000000000000000000000000",
13209 => "000000000000000000000000",
13210 => "000000000000000000000000",
13211 => "000000000000000000000000",
13212 => "000000000000000000000000",
13213 => "000000000000000000000000",
13214 => "000000000000000000000000",
13215 => "000000000000000000000000",
13216 => "000000000000000000000000",
13217 => "000000000000000000000000",
13218 => "000000000000000000000000",
13219 => "000000000000000000000000",
13220 => "000000000000000000000000",
13221 => "000000000000000000000000",
13222 => "000000000000000000000000",
13223 => "000000000000000000000000",
13224 => "000000000000000000000000",
13225 => "000000000000000000000000",
13226 => "000000000000000000000000",
13227 => "000000000000000000000000",
13228 => "000000000000000000000000",
13229 => "000000000000000000000000",
13230 => "000000000000000000000000",
13231 => "000000000000000000000000",
13232 => "000011010000110100001101",
13233 => "010000110100001101000011",
13234 => "010000110100001101000011",
13235 => "011000110110001101100011",
13236 => "011001100110011001100110",
13237 => "011001100110011001100110",
13238 => "011001100110011001100110",
13239 => "011000010110000101100001",
13240 => "010000110100001101000011",
13241 => "010000110100001101000011",
13242 => "010000110100001101000011",
13243 => "010000110100001101000011",
13244 => "010000110100001101000011",
13245 => "010000110100001101000011",
13246 => "010001110100011101000111",
13247 => "011001100110011001100110",
13248 => "011001100110011001100110",
13249 => "010010010100100101001001",
13250 => "010000110100001101000011",
13251 => "010000110100001101000011",
13252 => "010000110100001101000011",
13253 => "010000110100001101000011",
13254 => "010000110100001101000011",
13255 => "010000110100001101000011",
13256 => "010000110100001101000011",
13257 => "010000110100001101000011",
13258 => "010000110100001101000011",
13259 => "010000110100001101000011",
13260 => "010000110100001101000011",
13261 => "010000110100001101000011",
13262 => "010000110100001101000011",
13263 => "010000110100001101000011",
13264 => "010000110100001101000011",
13265 => "010000110100001101000011",
13266 => "010000110100001101000011",
13267 => "010000110100001101000011",
13268 => "010000110100001101000011",
13269 => "010000110100001101000011",
13270 => "010000110100001101000011",
13271 => "010000110100001101000011",
13272 => "010000110100001101000011",
13273 => "010000110100001101000011",
13274 => "010000110100001101000011",
13275 => "010000110100001101000011",
13276 => "010000110100001101000011",
13277 => "010000110100001101000011",
13278 => "010000110100001101000011",
13279 => "010000110100001101000011",
13280 => "010000110100001101000011",
13281 => "010000110100001101000011",
13282 => "010000110100001101000011",
13283 => "010000110100001101000011",
13284 => "010000110100001101000011",
13285 => "010000110100001101000011",
13286 => "010000110100001101000011",
13287 => "010000110100001101000011",
13288 => "010000110100001101000011",
13289 => "011001100110011001100110",
13290 => "011001100110011001100110",
13291 => "010100010101000101010001",
13292 => "010000110100001101000011",
13293 => "010000110100001101000011",
13294 => "010000110100001101000011",
13295 => "010000110100001101000011",
13296 => "010000110100001101000011",
13297 => "010000110100001101000011",
13298 => "010101110101011101010111",
13299 => "011001100110011001100110",
13300 => "011001100110011001100110",
13301 => "011001100110011001100110",
13302 => "011001100110011001100110",
13303 => "010001010100010101000101",
13304 => "010000110100001101000011",
13305 => "000111110001111100011111",
13306 => "000000000000000000000000",
13307 => "000000000000000000000000",
13308 => "000000000000000000000000",
13309 => "000000000000000000000000",
13310 => "000000000000000000000000",
13311 => "000000000000000000000000",
13312 => "000000000000000000000000",
13313 => "000000000000000000000000",
13314 => "000000000000000000000000",
13315 => "000000000000000000000000",
13316 => "000000000000000000000000",
13317 => "000000000000000000000000",
13318 => "000000000000000000000000",
13319 => "000000000000000000000000",
13320 => "000000000000000000000000",
13321 => "000000000000000000000000",
13322 => "000000000000000000000000",
13323 => "000000000000000000000000",
13324 => "000000000000000000000000",
13325 => "000000000000000000000000",
13326 => "000000000000000000000000",
13327 => "000000000000000000000000",
13328 => "000000000000000000000000",
13329 => "000000000000000000000000",
13330 => "000000000000000000000000",
13331 => "000000000000000000000000",
13332 => "000000000000000000000000",
13333 => "000000000000000000000000",
13334 => "000000000000000000000000",
13335 => "000000000000000000000000",
13336 => "000000000000000000000000",
13337 => "000000000000000000000000",
13338 => "000000000000000000000000",
13339 => "000000000000000000000000",
13340 => "000000000000000000000000",
13341 => "000000000000000000000000",
13342 => "000000000000000000000000",
13343 => "000000000000000000000000",
13344 => "000000000000000000000000",
13345 => "000000000000000000000000",
13346 => "000000000000000000000000",
13347 => "000000000000000000000000",
13348 => "000000000000000000000000",
13349 => "000000000000000000000000",
13350 => "000000000000000000000000",
13351 => "000000000000000000000000",
13352 => "000000000000000000000000",
13353 => "000000000000000000000000",
13354 => "000000000000000000000000",
13355 => "000000000000000000000000",
13356 => "000000000000000000000000",
13357 => "000000000000000000000000",
13358 => "000000000000000000000000",
13359 => "000000000000000000000000",
13360 => "000000000000000000000000",
13361 => "000000000000000000000000",
13362 => "000000000000000000000000",
13363 => "000000000000000000000000",
13364 => "000000000000000000000000",
13365 => "000000000000000000000000",
13366 => "000000000000000000000000",
13367 => "000000000000000000000000",
13368 => "000000000000000000000000",
13369 => "000000000000000000000000",
13370 => "000000000000000000000000",
13371 => "000000000000000000000000",
13372 => "000000000000000000000000",
13373 => "000000000000000000000000",
13374 => "000000000000000000000000",
13375 => "000000000000000000000000",
13376 => "000000000000000000000000",
13377 => "000000000000000000000000",
13378 => "001111110011111100111111",
13379 => "010000100100001001000010",
13380 => "010000100100001001000010",
13381 => "010000100100001001000010",
13382 => "010010010100100101001001",
13383 => "011001100110011001100110",
13384 => "011001100110011001100110",
13385 => "010001100100011001000110",
13386 => "010000110100001101000011",
13387 => "010000110100001101000011",
13388 => "010000110100001101000011",
13389 => "010000110100001101000011",
13390 => "010000110100001101000011",
13391 => "010000110100001101000011",
13392 => "010000110100001101000011",
13393 => "010000110100001101000011",
13394 => "010000110100001101000011",
13395 => "010000110100001101000011",
13396 => "010001110100011101000111",
13397 => "011001100110011001100110",
13398 => "011001100110011001100110",
13399 => "010010010100100101001001",
13400 => "010000110100001101000011",
13401 => "010000110100001101000011",
13402 => "010000110100001101000011",
13403 => "010000110100001101000011",
13404 => "010000110100001101000011",
13405 => "010000110100001101000011",
13406 => "010000110100001101000011",
13407 => "010000110100001101000011",
13408 => "010000110100001101000011",
13409 => "010000110100001101000011",
13410 => "010000110100001101000011",
13411 => "010000110100001101000011",
13412 => "010000110100001101000011",
13413 => "010000110100001101000011",
13414 => "010000110100001101000011",
13415 => "010000110100001101000011",
13416 => "010000110100001101000011",
13417 => "010000110100001101000011",
13418 => "010000110100001101000011",
13419 => "010000110100001101000011",
13420 => "010000110100001101000011",
13421 => "010000110100001101000011",
13422 => "010000110100001101000011",
13423 => "010000110100001101000011",
13424 => "010000110100001101000011",
13425 => "010000110100001101000011",
13426 => "010000110100001101000011",
13427 => "010000110100001101000011",
13428 => "010000110100001101000011",
13429 => "010000110100001101000011",
13430 => "010000110100001101000011",
13431 => "010000110100001101000011",
13432 => "010000110100001101000011",
13433 => "010000110100001101000011",
13434 => "010000110100001101000011",
13435 => "010000110100001101000011",
13436 => "010000110100001101000011",
13437 => "010000110100001101000011",
13438 => "010000110100001101000011",
13439 => "011001100110011001100110",
13440 => "011001100110011001100110",
13441 => "010100010101000101010001",
13442 => "010000110100001101000011",
13443 => "010000110100001101000011",
13444 => "010000110100001101000011",
13445 => "010000110100001101000011",
13446 => "010000110100001101000011",
13447 => "010000110100001101000011",
13448 => "010000110100001101000011",
13449 => "010000110100001101000011",
13450 => "010000110100001101000011",
13451 => "010000110100001101000011",
13452 => "010000110100001101000011",
13453 => "011001000110010001100100",
13454 => "011001100110011001100110",
13455 => "010100110101001101010011",
13456 => "010000100100001001000010",
13457 => "010000100100001001000010",
13458 => "010000100100001001000010",
13459 => "010000100100001001000010",
13460 => "000001100000011000000110",
13461 => "000000000000000000000000",
13462 => "000000000000000000000000",
13463 => "000000000000000000000000",
13464 => "000000000000000000000000",
13465 => "000000000000000000000000",
13466 => "000000000000000000000000",
13467 => "000000000000000000000000",
13468 => "000000000000000000000000",
13469 => "000000000000000000000000",
13470 => "000000000000000000000000",
13471 => "000000000000000000000000",
13472 => "000000000000000000000000",
13473 => "000000000000000000000000",
13474 => "000000000000000000000000",
13475 => "000000000000000000000000",
13476 => "000000000000000000000000",
13477 => "000000000000000000000000",
13478 => "000000000000000000000000",
13479 => "000000000000000000000000",
13480 => "000000000000000000000000",
13481 => "000000000000000000000000",
13482 => "000000000000000000000000",
13483 => "000000000000000000000000",
13484 => "000000000000000000000000",
13485 => "000000000000000000000000",
13486 => "000000000000000000000000",
13487 => "000000000000000000000000",
13488 => "000000000000000000000000",
13489 => "000000000000000000000000",
13490 => "000000000000000000000000",
13491 => "000000000000000000000000",
13492 => "000000000000000000000000",
13493 => "000000000000000000000000",
13494 => "000000000000000000000000",
13495 => "000000000000000000000000",
13496 => "000000000000000000000000",
13497 => "000000000000000000000000",
13498 => "000000000000000000000000",
13499 => "000000000000000000000000",
13500 => "000000000000000000000000",
13501 => "000000000000000000000000",
13502 => "000000000000000000000000",
13503 => "000000000000000000000000",
13504 => "000000000000000000000000",
13505 => "000000000000000000000000",
13506 => "000000000000000000000000",
13507 => "000000000000000000000000",
13508 => "000000000000000000000000",
13509 => "000000000000000000000000",
13510 => "000000000000000000000000",
13511 => "000000000000000000000000",
13512 => "000000000000000000000000",
13513 => "000000000000000000000000",
13514 => "000000000000000000000000",
13515 => "000000000000000000000000",
13516 => "000000000000000000000000",
13517 => "000000000000000000000000",
13518 => "000000000000000000000000",
13519 => "000000000000000000000000",
13520 => "000000000000000000000000",
13521 => "000000000000000000000000",
13522 => "000000000000000000000000",
13523 => "000000000000000000000000",
13524 => "000000000000000000000000",
13525 => "000000000000000000000000",
13526 => "000000000000000000000000",
13527 => "000000000000000000000000",
13528 => "001111110011111100111111",
13529 => "010000110100001101000011",
13530 => "010000110100001101000011",
13531 => "010000110100001101000011",
13532 => "010010100100101001001010",
13533 => "011001100110011001100110",
13534 => "011001100110011001100110",
13535 => "010001100100011001000110",
13536 => "010000110100001101000011",
13537 => "010000110100001101000011",
13538 => "010000110100001101000011",
13539 => "010000110100001101000011",
13540 => "010000110100001101000011",
13541 => "010000110100001101000011",
13542 => "010000110100001101000011",
13543 => "010000110100001101000011",
13544 => "010000110100001101000011",
13545 => "010000110100001101000011",
13546 => "010001110100011101000111",
13547 => "011001100110011001100110",
13548 => "011001100110011001100110",
13549 => "010010010100100101001001",
13550 => "010000110100001101000011",
13551 => "010000110100001101000011",
13552 => "010000110100001101000011",
13553 => "010000110100001101000011",
13554 => "010000110100001101000011",
13555 => "010000110100001101000011",
13556 => "010000110100001101000011",
13557 => "010000110100001101000011",
13558 => "010000110100001101000011",
13559 => "010000110100001101000011",
13560 => "010000110100001101000011",
13561 => "010000110100001101000011",
13562 => "010000110100001101000011",
13563 => "010000110100001101000011",
13564 => "010000110100001101000011",
13565 => "010000110100001101000011",
13566 => "010000110100001101000011",
13567 => "010000110100001101000011",
13568 => "010000110100001101000011",
13569 => "010000110100001101000011",
13570 => "010000110100001101000011",
13571 => "010000110100001101000011",
13572 => "010000110100001101000011",
13573 => "010000110100001101000011",
13574 => "010000110100001101000011",
13575 => "010000110100001101000011",
13576 => "010000110100001101000011",
13577 => "010000110100001101000011",
13578 => "010000110100001101000011",
13579 => "010000110100001101000011",
13580 => "010000110100001101000011",
13581 => "010000110100001101000011",
13582 => "010000110100001101000011",
13583 => "010000110100001101000011",
13584 => "010000110100001101000011",
13585 => "010000110100001101000011",
13586 => "010000110100001101000011",
13587 => "010000110100001101000011",
13588 => "010000110100001101000011",
13589 => "011001100110011001100110",
13590 => "011001100110011001100110",
13591 => "010100010101000101010001",
13592 => "010000110100001101000011",
13593 => "010000110100001101000011",
13594 => "010000110100001101000011",
13595 => "010000110100001101000011",
13596 => "010000110100001101000011",
13597 => "010000110100001101000011",
13598 => "010000110100001101000011",
13599 => "010000110100001101000011",
13600 => "010000110100001101000011",
13601 => "010000110100001101000011",
13602 => "010000110100001101000011",
13603 => "011001000110010001100100",
13604 => "011001100110011001100110",
13605 => "010100110101001101010011",
13606 => "010000110100001101000011",
13607 => "010000110100001101000011",
13608 => "010000110100001101000011",
13609 => "010000110100001101000011",
13610 => "000001100000011000000110",
13611 => "000000000000000000000000",
13612 => "000000000000000000000000",
13613 => "000000000000000000000000",
13614 => "000000000000000000000000",
13615 => "000000000000000000000000",
13616 => "000000000000000000000000",
13617 => "000000000000000000000000",
13618 => "000000000000000000000000",
13619 => "000000000000000000000000",
13620 => "000000000000000000000000",
13621 => "000000000000000000000000",
13622 => "000000000000000000000000",
13623 => "000000000000000000000000",
13624 => "000000000000000000000000",
13625 => "000000000000000000000000",
13626 => "000000000000000000000000",
13627 => "000000000000000000000000",
13628 => "000000000000000000000000",
13629 => "000000000000000000000000",
13630 => "000000000000000000000000",
13631 => "000000000000000000000000",
13632 => "000000000000000000000000",
13633 => "000000000000000000000000",
13634 => "000000000000000000000000",
13635 => "000000000000000000000000",
13636 => "000000000000000000000000",
13637 => "000000000000000000000000",
13638 => "000000000000000000000000",
13639 => "000000000000000000000000",
13640 => "000000000000000000000000",
13641 => "000000000000000000000000",
13642 => "000000000000000000000000",
13643 => "000000000000000000000000",
13644 => "000000000000000000000000",
13645 => "000000000000000000000000",
13646 => "000000000000000000000000",
13647 => "000000000000000000000000",
13648 => "000000000000000000000000",
13649 => "000000000000000000000000",
13650 => "000000000000000000000000",
13651 => "000000000000000000000000",
13652 => "000000000000000000000000",
13653 => "000000000000000000000000",
13654 => "000000000000000000000000",
13655 => "000000000000000000000000",
13656 => "000000000000000000000000",
13657 => "000000000000000000000000",
13658 => "000000000000000000000000",
13659 => "000000000000000000000000",
13660 => "000000000000000000000000",
13661 => "000000000000000000000000",
13662 => "000000000000000000000000",
13663 => "000000000000000000000000",
13664 => "000000000000000000000000",
13665 => "000000000000000000000000",
13666 => "000000000000000000000000",
13667 => "000000000000000000000000",
13668 => "000000000000000000000000",
13669 => "000000000000000000000000",
13670 => "000000000000000000000000",
13671 => "000000000000000000000000",
13672 => "000000000000000000000000",
13673 => "000000000000000000000000",
13674 => "000000000000000000000000",
13675 => "000010010000100100001001",
13676 => "001010000010100000101000",
13677 => "001010000010100000101000",
13678 => "010101010101010101010101",
13679 => "010110000101100001011000",
13680 => "010110000101100001011000",
13681 => "010110000101100001011000",
13682 => "010101110101011101010111",
13683 => "010100010101000101010001",
13684 => "010100010101000101010001",
13685 => "010001000100010001000100",
13686 => "010000110100001101000011",
13687 => "010000110100001101000011",
13688 => "010000110100001101000011",
13689 => "010001100100011001000110",
13690 => "010110000101100001011000",
13691 => "010110000101100001011000",
13692 => "010001010100010101000101",
13693 => "010000110100001101000011",
13694 => "010000110100001101000011",
13695 => "010000110100001101000011",
13696 => "010001110100011101000111",
13697 => "011001100110011001100110",
13698 => "011001100110011001100110",
13699 => "010010010100100101001001",
13700 => "010000110100001101000011",
13701 => "010000110100001101000011",
13702 => "010000110100001101000011",
13703 => "010000110100001101000011",
13704 => "010000110100001101000011",
13705 => "010000110100001101000011",
13706 => "010000110100001101000011",
13707 => "010000110100001101000011",
13708 => "010000110100001101000011",
13709 => "010000110100001101000011",
13710 => "010000110100001101000011",
13711 => "010000110100001101000011",
13712 => "010000110100001101000011",
13713 => "010000110100001101000011",
13714 => "010000110100001101000011",
13715 => "010000110100001101000011",
13716 => "010000110100001101000011",
13717 => "010000110100001101000011",
13718 => "010000110100001101000011",
13719 => "010000110100001101000011",
13720 => "010000110100001101000011",
13721 => "010000110100001101000011",
13722 => "010000110100001101000011",
13723 => "010000110100001101000011",
13724 => "010000110100001101000011",
13725 => "010000110100001101000011",
13726 => "010000110100001101000011",
13727 => "010000110100001101000011",
13728 => "010000110100001101000011",
13729 => "010000110100001101000011",
13730 => "010000110100001101000011",
13731 => "010000110100001101000011",
13732 => "010000110100001101000011",
13733 => "010000110100001101000011",
13734 => "010000110100001101000011",
13735 => "010000110100001101000011",
13736 => "010000110100001101000011",
13737 => "010000110100001101000011",
13738 => "010000110100001101000011",
13739 => "011001100110011001100110",
13740 => "011001100110011001100110",
13741 => "010100010101000101010001",
13742 => "010000110100001101000011",
13743 => "010000110100001101000011",
13744 => "010000110100001101000011",
13745 => "010000110100001101000011",
13746 => "010101110101011101010111",
13747 => "010110000101100001011000",
13748 => "010011000100110001001100",
13749 => "010000110100001101000011",
13750 => "010000110100001101000011",
13751 => "010000110100001101000011",
13752 => "010000110100001101000011",
13753 => "010100000101000001010000",
13754 => "010100010101000101010001",
13755 => "010101010101010101010101",
13756 => "010110000101100001011000",
13757 => "010110000101100001011000",
13758 => "010110000101100001011000",
13759 => "010110000101100001011000",
13760 => "001011000010110000101100",
13761 => "001010000010100000101000",
13762 => "000101000001010000010100",
13763 => "000000000000000000000000",
13764 => "000000000000000000000000",
13765 => "000000000000000000000000",
13766 => "000000000000000000000000",
13767 => "000000000000000000000000",
13768 => "000000000000000000000000",
13769 => "000000000000000000000000",
13770 => "000000000000000000000000",
13771 => "000000000000000000000000",
13772 => "000000000000000000000000",
13773 => "000000000000000000000000",
13774 => "000000000000000000000000",
13775 => "000000000000000000000000",
13776 => "000000000000000000000000",
13777 => "000000000000000000000000",
13778 => "000000000000000000000000",
13779 => "000000000000000000000000",
13780 => "000000000000000000000000",
13781 => "000000000000000000000000",
13782 => "000000000000000000000000",
13783 => "000000000000000000000000",
13784 => "000000000000000000000000",
13785 => "000000000000000000000000",
13786 => "000000000000000000000000",
13787 => "000000000000000000000000",
13788 => "000000000000000000000000",
13789 => "000000000000000000000000",
13790 => "000000000000000000000000",
13791 => "000000000000000000000000",
13792 => "000000000000000000000000",
13793 => "000000000000000000000000",
13794 => "000000000000000000000000",
13795 => "000000000000000000000000",
13796 => "000000000000000000000000",
13797 => "000000000000000000000000",
13798 => "000000000000000000000000",
13799 => "000000000000000000000000",
13800 => "000000000000000000000000",
13801 => "000000000000000000000000",
13802 => "000000000000000000000000",
13803 => "000000000000000000000000",
13804 => "000000000000000000000000",
13805 => "000000000000000000000000",
13806 => "000000000000000000000000",
13807 => "000000000000000000000000",
13808 => "000000000000000000000000",
13809 => "000000000000000000000000",
13810 => "000000000000000000000000",
13811 => "000000000000000000000000",
13812 => "000000000000000000000000",
13813 => "000000000000000000000000",
13814 => "000000000000000000000000",
13815 => "000000000000000000000000",
13816 => "000000000000000000000000",
13817 => "000000000000000000000000",
13818 => "000000000000000000000000",
13819 => "000000000000000000000000",
13820 => "000000000000000000000000",
13821 => "000000000000000000000000",
13822 => "000000000000000000000000",
13823 => "000000000000000000000000",
13824 => "000000000000000000000000",
13825 => "000011110000111100001111",
13826 => "010000110100001101000011",
13827 => "010000110100001101000011",
13828 => "011001000110010001100100",
13829 => "011001100110011001100110",
13830 => "011001100110011001100110",
13831 => "011001100110011001100110",
13832 => "010111110101111101011111",
13833 => "010000110100001101000011",
13834 => "010000110100001101000011",
13835 => "010000110100001101000011",
13836 => "010000110100001101000011",
13837 => "010000110100001101000011",
13838 => "010000110100001101000011",
13839 => "010010000100100001001000",
13840 => "011001100110011001100110",
13841 => "011001100110011001100110",
13842 => "010001110100011101000111",
13843 => "010000110100001101000011",
13844 => "010000110100001101000011",
13845 => "010000110100001101000011",
13846 => "010001110100011101000111",
13847 => "011001100110011001100110",
13848 => "011001100110011001100110",
13849 => "010010010100100101001001",
13850 => "010000110100001101000011",
13851 => "010000110100001101000011",
13852 => "010000110100001101000011",
13853 => "010000110100001101000011",
13854 => "010000110100001101000011",
13855 => "010000110100001101000011",
13856 => "010000110100001101000011",
13857 => "010000110100001101000011",
13858 => "010000110100001101000011",
13859 => "010000110100001101000011",
13860 => "010000110100001101000011",
13861 => "010000110100001101000011",
13862 => "010000110100001101000011",
13863 => "010000110100001101000011",
13864 => "010000110100001101000011",
13865 => "010000110100001101000011",
13866 => "010000110100001101000011",
13867 => "010000110100001101000011",
13868 => "010000110100001101000011",
13869 => "010000110100001101000011",
13870 => "010000110100001101000011",
13871 => "010000110100001101000011",
13872 => "010000110100001101000011",
13873 => "010000110100001101000011",
13874 => "010000110100001101000011",
13875 => "010000110100001101000011",
13876 => "010000110100001101000011",
13877 => "010000110100001101000011",
13878 => "010000110100001101000011",
13879 => "010000110100001101000011",
13880 => "010000110100001101000011",
13881 => "010000110100001101000011",
13882 => "010000110100001101000011",
13883 => "010000110100001101000011",
13884 => "010000110100001101000011",
13885 => "010000110100001101000011",
13886 => "010000110100001101000011",
13887 => "010000110100001101000011",
13888 => "010000110100001101000011",
13889 => "011001100110011001100110",
13890 => "011001100110011001100110",
13891 => "010100010101000101010001",
13892 => "010000110100001101000011",
13893 => "010000110100001101000011",
13894 => "010000110100001101000011",
13895 => "010000110100001101000011",
13896 => "011001010110010101100101",
13897 => "011001100110011001100110",
13898 => "010100100101001001010010",
13899 => "010000110100001101000011",
13900 => "010000110100001101000011",
13901 => "010000110100001101000011",
13902 => "010000110100001101000011",
13903 => "010000110100001101000011",
13904 => "010000110100001101000011",
13905 => "010101100101011001010110",
13906 => "011001100110011001100110",
13907 => "011001100110011001100110",
13908 => "011001100110011001100110",
13909 => "011001100110011001100110",
13910 => "010001100100011001000110",
13911 => "010000110100001101000011",
13912 => "001000100010001000100010",
13913 => "000000000000000000000000",
13914 => "000000000000000000000000",
13915 => "000000000000000000000000",
13916 => "000000000000000000000000",
13917 => "000000000000000000000000",
13918 => "000000000000000000000000",
13919 => "000000000000000000000000",
13920 => "000000000000000000000000",
13921 => "000000000000000000000000",
13922 => "000000000000000000000000",
13923 => "000000000000000000000000",
13924 => "000000000000000000000000",
13925 => "000000000000000000000000",
13926 => "000000000000000000000000",
13927 => "000000000000000000000000",
13928 => "000000000000000000000000",
13929 => "000000000000000000000000",
13930 => "000000000000000000000000",
13931 => "000000000000000000000000",
13932 => "000000000000000000000000",
13933 => "000000000000000000000000",
13934 => "000000000000000000000000",
13935 => "000000000000000000000000",
13936 => "000000000000000000000000",
13937 => "000000000000000000000000",
13938 => "000000000000000000000000",
13939 => "000000000000000000000000",
13940 => "000000000000000000000000",
13941 => "000000000000000000000000",
13942 => "000000000000000000000000",
13943 => "000000000000000000000000",
13944 => "000000000000000000000000",
13945 => "000000000000000000000000",
13946 => "000000000000000000000000",
13947 => "000000000000000000000000",
13948 => "000000000000000000000000",
13949 => "000000000000000000000000",
13950 => "000000000000000000000000",
13951 => "000000000000000000000000",
13952 => "000000000000000000000000",
13953 => "000000000000000000000000",
13954 => "000000000000000000000000",
13955 => "000000000000000000000000",
13956 => "000000000000000000000000",
13957 => "000000000000000000000000",
13958 => "000000000000000000000000",
13959 => "000000000000000000000000",
13960 => "000000000000000000000000",
13961 => "000000000000000000000000",
13962 => "000000000000000000000000",
13963 => "000000000000000000000000",
13964 => "000000000000000000000000",
13965 => "000000000000000000000000",
13966 => "000000000000000000000000",
13967 => "000000000000000000000000",
13968 => "000000000000000000000000",
13969 => "000000000000000000000000",
13970 => "000000000000000000000000",
13971 => "000100000001000000010000",
13972 => "000100010001000100010001",
13973 => "000101100001011000010110",
13974 => "000110100001101000011010",
13975 => "001001000010010000100100",
13976 => "010011000100110001001100",
13977 => "010011000100110001001100",
13978 => "010111000101110001011100",
13979 => "010111010101110101011101",
13980 => "010111010101110101011101",
13981 => "010111010101110101011101",
13982 => "010110000101100001011000",
13983 => "010000110100001101000011",
13984 => "010000110100001101000011",
13985 => "010000110100001101000011",
13986 => "010000110100001101000011",
13987 => "010000110100001101000011",
13988 => "010000110100001101000011",
13989 => "010010000100100001001000",
13990 => "011001100110011001100110",
13991 => "011001100110011001100110",
13992 => "010001110100011101000111",
13993 => "010000110100001101000011",
13994 => "010000110100001101000011",
13995 => "010000110100001101000011",
13996 => "010001110100011101000111",
13997 => "011001100110011001100110",
13998 => "011001100110011001100110",
13999 => "010010010100100101001001",
14000 => "010000110100001101000011",
14001 => "010000110100001101000011",
14002 => "010000110100001101000011",
14003 => "010000110100001101000011",
14004 => "010000110100001101000011",
14005 => "010000110100001101000011",
14006 => "010000110100001101000011",
14007 => "010000110100001101000011",
14008 => "010000110100001101000011",
14009 => "010000110100001101000011",
14010 => "010001000100010001000100",
14011 => "010011000100110001001100",
14012 => "010011000100110001001100",
14013 => "010001010100010101000101",
14014 => "010000110100001101000011",
14015 => "010000110100001101000011",
14016 => "010000110100001101000011",
14017 => "010000110100001101000011",
14018 => "010000110100001101000011",
14019 => "010000110100001101000011",
14020 => "010000110100001101000011",
14021 => "010000110100001101000011",
14022 => "010000110100001101000011",
14023 => "010000110100001101000011",
14024 => "010000110100001101000011",
14025 => "010011000100110001001100",
14026 => "010011000100110001001100",
14027 => "010001100100011001000110",
14028 => "010000110100001101000011",
14029 => "010000110100001101000011",
14030 => "010000110100001101000011",
14031 => "010000110100001101000011",
14032 => "010000110100001101000011",
14033 => "010000110100001101000011",
14034 => "010000110100001101000011",
14035 => "010000110100001101000011",
14036 => "010000110100001101000011",
14037 => "010000110100001101000011",
14038 => "010000110100001101000011",
14039 => "011001100110011001100110",
14040 => "011001100110011001100110",
14041 => "010100010101000101010001",
14042 => "010000110100001101000011",
14043 => "010000110100001101000011",
14044 => "010000110100001101000011",
14045 => "010000110100001101000011",
14046 => "011001010110010101100101",
14047 => "011001100110011001100110",
14048 => "010100100101001001010010",
14049 => "010000110100001101000011",
14050 => "010000110100001101000011",
14051 => "010000110100001101000011",
14052 => "010000110100001101000011",
14053 => "010000110100001101000011",
14054 => "010000110100001101000011",
14055 => "010100010101000101010001",
14056 => "010111010101110101011101",
14057 => "010111010101110101011101",
14058 => "010111010101110101011101",
14059 => "010111010101110101011101",
14060 => "010011010100110101001101",
14061 => "010011000100110001001100",
14062 => "001100110011001100110011",
14063 => "000110100001101000011010",
14064 => "000110000001100000011000",
14065 => "000100010001000100010001",
14066 => "000100010001000100010001",
14067 => "000000100000001000000010",
14068 => "000000000000000000000000",
14069 => "000000000000000000000000",
14070 => "000000000000000000000000",
14071 => "000000000000000000000000",
14072 => "000000000000000000000000",
14073 => "000000000000000000000000",
14074 => "000000000000000000000000",
14075 => "000000000000000000000000",
14076 => "000000000000000000000000",
14077 => "000000000000000000000000",
14078 => "000000000000000000000000",
14079 => "000000000000000000000000",
14080 => "000000000000000000000000",
14081 => "000000000000000000000000",
14082 => "000000000000000000000000",
14083 => "000000000000000000000000",
14084 => "000000000000000000000000",
14085 => "000000000000000000000000",
14086 => "000000000000000000000000",
14087 => "000000000000000000000000",
14088 => "000000000000000000000000",
14089 => "000000000000000000000000",
14090 => "000000000000000000000000",
14091 => "000000000000000000000000",
14092 => "000000000000000000000000",
14093 => "000000000000000000000000",
14094 => "000000000000000000000000",
14095 => "000000000000000000000000",
14096 => "000000000000000000000000",
14097 => "000000000000000000000000",
14098 => "000000000000000000000000",
14099 => "000000000000000000000000",
14100 => "000000000000000000000000",
14101 => "000000000000000000000000",
14102 => "000000000000000000000000",
14103 => "000000000000000000000000",
14104 => "000000000000000000000000",
14105 => "000000000000000000000000",
14106 => "000000000000000000000000",
14107 => "000000000000000000000000",
14108 => "000000000000000000000000",
14109 => "000000000000000000000000",
14110 => "000000000000000000000000",
14111 => "000000000000000000000000",
14112 => "000000000000000000000000",
14113 => "000000000000000000000000",
14114 => "000000000000000000000000",
14115 => "000000000000000000000000",
14116 => "000000000000000000000000",
14117 => "000000000000000000000000",
14118 => "000000000000000000000000",
14119 => "000000000000000000000000",
14120 => "000000000000000000000000",
14121 => "010000010100000101000001",
14122 => "010000110100001101000011",
14123 => "010101110101011101010111",
14124 => "011001100110011001100110",
14125 => "011001100110011001100110",
14126 => "011001100110011001100110",
14127 => "011001100110011001100110",
14128 => "010001010100010101000101",
14129 => "010000110100001101000011",
14130 => "010000110100001101000011",
14131 => "010000110100001101000011",
14132 => "010000110100001101000011",
14133 => "010000110100001101000011",
14134 => "010000110100001101000011",
14135 => "010000110100001101000011",
14136 => "010000110100001101000011",
14137 => "010000110100001101000011",
14138 => "010000110100001101000011",
14139 => "010010000100100001001000",
14140 => "011001100110011001100110",
14141 => "011001100110011001100110",
14142 => "010001110100011101000111",
14143 => "010000110100001101000011",
14144 => "010000110100001101000011",
14145 => "010000110100001101000011",
14146 => "010001110100011101000111",
14147 => "011001100110011001100110",
14148 => "011001100110011001100110",
14149 => "010010010100100101001001",
14150 => "010000110100001101000011",
14151 => "010000110100001101000011",
14152 => "010000110100001101000011",
14153 => "010000110100001101000011",
14154 => "010000110100001101000011",
14155 => "010000110100001101000011",
14156 => "010000110100001101000011",
14157 => "010000110100001101000011",
14158 => "010000110100001101000011",
14159 => "010000110100001101000011",
14160 => "010001010100010101000101",
14161 => "011001100110011001100110",
14162 => "011001100110011001100110",
14163 => "010011000100110001001100",
14164 => "010000110100001101000011",
14165 => "010000110100001101000011",
14166 => "010000110100001101000011",
14167 => "010000110100001101000011",
14168 => "010000110100001101000011",
14169 => "010000110100001101000011",
14170 => "010000110100001101000011",
14171 => "010000110100001101000011",
14172 => "010000110100001101000011",
14173 => "010000110100001101000011",
14174 => "010000110100001101000011",
14175 => "011001100110011001100110",
14176 => "011001100110011001100110",
14177 => "010011110100111101001111",
14178 => "010000110100001101000011",
14179 => "010000110100001101000011",
14180 => "010000110100001101000011",
14181 => "010000110100001101000011",
14182 => "010000110100001101000011",
14183 => "010000110100001101000011",
14184 => "010000110100001101000011",
14185 => "010000110100001101000011",
14186 => "010000110100001101000011",
14187 => "010000110100001101000011",
14188 => "010000110100001101000011",
14189 => "011001100110011001100110",
14190 => "011001100110011001100110",
14191 => "010100010101000101010001",
14192 => "010000110100001101000011",
14193 => "010000110100001101000011",
14194 => "010000110100001101000011",
14195 => "010000110100001101000011",
14196 => "011001010110010101100101",
14197 => "011001100110011001100110",
14198 => "010100100101001001010010",
14199 => "010000110100001101000011",
14200 => "010000110100001101000011",
14201 => "010000110100001101000011",
14202 => "010000110100001101000011",
14203 => "010000110100001101000011",
14204 => "010000110100001101000011",
14205 => "010000110100001101000011",
14206 => "010000110100001101000011",
14207 => "010000110100001101000011",
14208 => "010000110100001101000011",
14209 => "010000110100001101000011",
14210 => "011000110110001101100011",
14211 => "011001100110011001100110",
14212 => "011001100110011001100110",
14213 => "011001100110011001100110",
14214 => "011000010110000101100001",
14215 => "010000110100001101000011",
14216 => "010000110100001101000011",
14217 => "000010000000100000001000",
14218 => "000000000000000000000000",
14219 => "000000000000000000000000",
14220 => "000000000000000000000000",
14221 => "000000000000000000000000",
14222 => "000000000000000000000000",
14223 => "000000000000000000000000",
14224 => "000000000000000000000000",
14225 => "000000000000000000000000",
14226 => "000000000000000000000000",
14227 => "000000000000000000000000",
14228 => "000000000000000000000000",
14229 => "000000000000000000000000",
14230 => "000000000000000000000000",
14231 => "000000000000000000000000",
14232 => "000000000000000000000000",
14233 => "000000000000000000000000",
14234 => "000000000000000000000000",
14235 => "000000000000000000000000",
14236 => "000000000000000000000000",
14237 => "000000000000000000000000",
14238 => "000000000000000000000000",
14239 => "000000000000000000000000",
14240 => "000000000000000000000000",
14241 => "000000000000000000000000",
14242 => "000000000000000000000000",
14243 => "000000000000000000000000",
14244 => "000000000000000000000000",
14245 => "000000000000000000000000",
14246 => "000000000000000000000000",
14247 => "000000000000000000000000",
14248 => "000000000000000000000000",
14249 => "000000000000000000000000",
14250 => "000000000000000000000000",
14251 => "000000000000000000000000",
14252 => "000000000000000000000000",
14253 => "000000000000000000000000",
14254 => "000000000000000000000000",
14255 => "000000000000000000000000",
14256 => "000000000000000000000000",
14257 => "000000000000000000000000",
14258 => "000000000000000000000000",
14259 => "000000000000000000000000",
14260 => "000000000000000000000000",
14261 => "000000000000000000000000",
14262 => "000000000000000000000000",
14263 => "000000000000000000000000",
14264 => "000000000000000000000000",
14265 => "000000000000000000000000",
14266 => "000000000000000000000000",
14267 => "000000000000000000000000",
14268 => "000000000000000000000000",
14269 => "000000000000000000000000",
14270 => "000000000000000000000000",
14271 => "010000010100000101000001",
14272 => "010000110100001101000011",
14273 => "010101110101011101010111",
14274 => "011001100110011001100110",
14275 => "011001100110011001100110",
14276 => "011001100110011001100110",
14277 => "011001100110011001100110",
14278 => "010001010100010101000101",
14279 => "010000110100001101000011",
14280 => "010000110100001101000011",
14281 => "010000110100001101000011",
14282 => "010000110100001101000011",
14283 => "010000110100001101000011",
14284 => "010000110100001101000011",
14285 => "010000110100001101000011",
14286 => "010000110100001101000011",
14287 => "010000110100001101000011",
14288 => "010000110100001101000011",
14289 => "010010000100100001001000",
14290 => "011001100110011001100110",
14291 => "011001100110011001100110",
14292 => "010001110100011101000111",
14293 => "010000110100001101000011",
14294 => "010000110100001101000011",
14295 => "010000110100001101000011",
14296 => "010001110100011101000111",
14297 => "011001100110011001100110",
14298 => "011001100110011001100110",
14299 => "010010010100100101001001",
14300 => "010000110100001101000011",
14301 => "010000110100001101000011",
14302 => "010000110100001101000011",
14303 => "010000110100001101000011",
14304 => "010000110100001101000011",
14305 => "010000110100001101000011",
14306 => "010000110100001101000011",
14307 => "010000110100001101000011",
14308 => "010000110100001101000011",
14309 => "010000110100001101000011",
14310 => "010001010100010101000101",
14311 => "011001100110011001100110",
14312 => "011001100110011001100110",
14313 => "010011000100110001001100",
14314 => "010000110100001101000011",
14315 => "010000110100001101000011",
14316 => "010000110100001101000011",
14317 => "010000110100001101000011",
14318 => "010000110100001101000011",
14319 => "010000110100001101000011",
14320 => "010000110100001101000011",
14321 => "010000110100001101000011",
14322 => "010000110100001101000011",
14323 => "010000110100001101000011",
14324 => "010000110100001101000011",
14325 => "011001100110011001100110",
14326 => "011001100110011001100110",
14327 => "010011110100111101001111",
14328 => "010000110100001101000011",
14329 => "010000110100001101000011",
14330 => "010000110100001101000011",
14331 => "010000110100001101000011",
14332 => "010000110100001101000011",
14333 => "010000110100001101000011",
14334 => "010000110100001101000011",
14335 => "010000110100001101000011",
14336 => "010000110100001101000011",
14337 => "010000110100001101000011",
14338 => "010000110100001101000011",
14339 => "011001100110011001100110",
14340 => "011001100110011001100110",
14341 => "010100010101000101010001",
14342 => "010000110100001101000011",
14343 => "010000110100001101000011",
14344 => "010000110100001101000011",
14345 => "010000110100001101000011",
14346 => "011001010110010101100101",
14347 => "011001100110011001100110",
14348 => "010100100101001001010010",
14349 => "010000110100001101000011",
14350 => "010000110100001101000011",
14351 => "010000110100001101000011",
14352 => "010000110100001101000011",
14353 => "010000110100001101000011",
14354 => "010000110100001101000011",
14355 => "010000110100001101000011",
14356 => "010000110100001101000011",
14357 => "010000110100001101000011",
14358 => "010000110100001101000011",
14359 => "010000110100001101000011",
14360 => "011000110110001101100011",
14361 => "011001100110011001100110",
14362 => "011001100110011001100110",
14363 => "011001100110011001100110",
14364 => "011000010110000101100001",
14365 => "010000110100001101000011",
14366 => "010000110100001101000011",
14367 => "000010000000100000001000",
14368 => "000000000000000000000000",
14369 => "000000000000000000000000",
14370 => "000000000000000000000000",
14371 => "000000000000000000000000",
14372 => "000000000000000000000000",
14373 => "000000000000000000000000",
14374 => "000000000000000000000000",
14375 => "000000000000000000000000",
14376 => "000000000000000000000000",
14377 => "000000000000000000000000",
14378 => "000000000000000000000000",
14379 => "000000000000000000000000",
14380 => "000000000000000000000000",
14381 => "000000000000000000000000",
14382 => "000000000000000000000000",
14383 => "000000000000000000000000",
14384 => "000000000000000000000000",
14385 => "000000000000000000000000",
14386 => "000000000000000000000000",
14387 => "000000000000000000000000",
14388 => "000000000000000000000000",
14389 => "000000000000000000000000",
14390 => "000000000000000000000000",
14391 => "000000000000000000000000",
14392 => "000000000000000000000000",
14393 => "000000000000000000000000",
14394 => "000000000000000000000000",
14395 => "000000000000000000000000",
14396 => "000000000000000000000000",
14397 => "000000000000000000000000",
14398 => "000000000000000000000000",
14399 => "000000000000000000000000",
14400 => "000000000000000000000000",
14401 => "000000000000000000000000",
14402 => "000000000000000000000000",
14403 => "000000000000000000000000",
14404 => "000000000000000000000000",
14405 => "000000000000000000000000",
14406 => "000000000000000000000000",
14407 => "000000000000000000000000",
14408 => "000000000000000000000000",
14409 => "000000000000000000000000",
14410 => "000000000000000000000000",
14411 => "000000000000000000000000",
14412 => "000000000000000000000000",
14413 => "000000000000000000000000",
14414 => "000000000000000000000000",
14415 => "000000000000000000000000",
14416 => "001001110010011100100111",
14417 => "010000010100000101000001",
14418 => "010000010100000101000001",
14419 => "010000010100000101000001",
14420 => "010000010100000101000001",
14421 => "010000110100001101000011",
14422 => "010000110100001101000011",
14423 => "010001000100010001000100",
14424 => "010001000100010001000100",
14425 => "010001000100010001000100",
14426 => "010001000100010001000100",
14427 => "010001000100010001000100",
14428 => "010000110100001101000011",
14429 => "010000110100001101000011",
14430 => "010000110100001101000011",
14431 => "010000110100001101000011",
14432 => "010000110100001101000011",
14433 => "010000110100001101000011",
14434 => "010000110100001101000011",
14435 => "010000110100001101000011",
14436 => "010000110100001101000011",
14437 => "010000110100001101000011",
14438 => "010000110100001101000011",
14439 => "010010000100100001001000",
14440 => "011001100110011001100110",
14441 => "011001100110011001100110",
14442 => "010001110100011101000111",
14443 => "010000110100001101000011",
14444 => "010000110100001101000011",
14445 => "010000110100001101000011",
14446 => "010001110100011101000111",
14447 => "011001100110011001100110",
14448 => "011001100110011001100110",
14449 => "010010010100100101001001",
14450 => "010000110100001101000011",
14451 => "010000110100001101000011",
14452 => "010000110100001101000011",
14453 => "010000110100001101000011",
14454 => "010000110100001101000011",
14455 => "010000110100001101000011",
14456 => "010000110100001101000011",
14457 => "010000110100001101000011",
14458 => "010100010101000101010001",
14459 => "011001010110010101100101",
14460 => "011000110110001101100011",
14461 => "010001000100010001000100",
14462 => "010001000100010001000100",
14463 => "010111000101110001011100",
14464 => "011001010110010101100101",
14465 => "010110000101100001011000",
14466 => "010000110100001101000011",
14467 => "010000110100001101000011",
14468 => "010000110100001101000011",
14469 => "010000110100001101000011",
14470 => "010000110100001101000011",
14471 => "010000110100001101000011",
14472 => "010011110100111101001111",
14473 => "011001010110010101100101",
14474 => "011001010110010101100101",
14475 => "010001000100010001000100",
14476 => "010001000100010001000100",
14477 => "010110100101101001011010",
14478 => "011001010110010101100101",
14479 => "010110100101101001011010",
14480 => "010000110100001101000011",
14481 => "010000110100001101000011",
14482 => "010000110100001101000011",
14483 => "010000110100001101000011",
14484 => "010000110100001101000011",
14485 => "010000110100001101000011",
14486 => "010000110100001101000011",
14487 => "010000110100001101000011",
14488 => "010000110100001101000011",
14489 => "011001100110011001100110",
14490 => "011001100110011001100110",
14491 => "010100010101000101010001",
14492 => "010000110100001101000011",
14493 => "010000110100001101000011",
14494 => "010000110100001101000011",
14495 => "010000110100001101000011",
14496 => "011001010110010101100101",
14497 => "011001100110011001100110",
14498 => "010100100101001001010010",
14499 => "010000110100001101000011",
14500 => "010000110100001101000011",
14501 => "010000110100001101000011",
14502 => "010000110100001101000011",
14503 => "010000110100001101000011",
14504 => "010000110100001101000011",
14505 => "010000110100001101000011",
14506 => "010000110100001101000011",
14507 => "010000110100001101000011",
14508 => "010000110100001101000011",
14509 => "010000110100001101000011",
14510 => "010001000100010001000100",
14511 => "010001000100010001000100",
14512 => "010001000100010001000100",
14513 => "010001000100010001000100",
14514 => "010001000100010001000100",
14515 => "010000110100001101000011",
14516 => "010000110100001101000011",
14517 => "010000010100000101000001",
14518 => "010000010100000101000001",
14519 => "010000010100000101000001",
14520 => "010000010100000101000001",
14521 => "001110010011100100111001",
14522 => "000000000000000000000000",
14523 => "000000000000000000000000",
14524 => "000000000000000000000000",
14525 => "000000000000000000000000",
14526 => "000000000000000000000000",
14527 => "000000000000000000000000",
14528 => "000000000000000000000000",
14529 => "000000000000000000000000",
14530 => "000000000000000000000000",
14531 => "000000000000000000000000",
14532 => "000000000000000000000000",
14533 => "000000000000000000000000",
14534 => "000000000000000000000000",
14535 => "000000000000000000000000",
14536 => "000000000000000000000000",
14537 => "000000000000000000000000",
14538 => "000000000000000000000000",
14539 => "000000000000000000000000",
14540 => "000000000000000000000000",
14541 => "000000000000000000000000",
14542 => "000000000000000000000000",
14543 => "000000000000000000000000",
14544 => "000000000000000000000000",
14545 => "000000000000000000000000",
14546 => "000000000000000000000000",
14547 => "000000000000000000000000",
14548 => "000000000000000000000000",
14549 => "000000000000000000000000",
14550 => "000000000000000000000000",
14551 => "000000000000000000000000",
14552 => "000000000000000000000000",
14553 => "000000000000000000000000",
14554 => "000000000000000000000000",
14555 => "000000000000000000000000",
14556 => "000000000000000000000000",
14557 => "000000000000000000000000",
14558 => "000000000000000000000000",
14559 => "000000000000000000000000",
14560 => "000000000000000000000000",
14561 => "000000000000000000000000",
14562 => "000000000000000000000000",
14563 => "000000000000000000000000",
14564 => "000000000000000000000000",
14565 => "000000000000000000000000",
14566 => "001010000010100000101000",
14567 => "010000110100001101000011",
14568 => "010000110100001101000011",
14569 => "010000110100001101000011",
14570 => "010000110100001101000011",
14571 => "010000110100001101000011",
14572 => "010000110100001101000011",
14573 => "010000110100001101000011",
14574 => "010000110100001101000011",
14575 => "010000110100001101000011",
14576 => "010000110100001101000011",
14577 => "010000110100001101000011",
14578 => "010000110100001101000011",
14579 => "010000110100001101000011",
14580 => "010000110100001101000011",
14581 => "010000110100001101000011",
14582 => "010000110100001101000011",
14583 => "010000110100001101000011",
14584 => "010000110100001101000011",
14585 => "010000110100001101000011",
14586 => "010000110100001101000011",
14587 => "010000110100001101000011",
14588 => "010000110100001101000011",
14589 => "010010000100100001001000",
14590 => "011001100110011001100110",
14591 => "011001100110011001100110",
14592 => "010001110100011101000111",
14593 => "010000110100001101000011",
14594 => "010000110100001101000011",
14595 => "010000110100001101000011",
14596 => "010001110100011101000111",
14597 => "011001100110011001100110",
14598 => "011001100110011001100110",
14599 => "010010010100100101001001",
14600 => "010000110100001101000011",
14601 => "010000110100001101000011",
14602 => "010000110100001101000011",
14603 => "010000110100001101000011",
14604 => "010000110100001101000011",
14605 => "010000110100001101000011",
14606 => "010000110100001101000011",
14607 => "010000110100001101000011",
14608 => "010100010101000101010001",
14609 => "011001100110011001100110",
14610 => "011001000110010001100100",
14611 => "010000110100001101000011",
14612 => "010000110100001101000011",
14613 => "010111010101110101011101",
14614 => "011001100110011001100110",
14615 => "010110010101100101011001",
14616 => "010000110100001101000011",
14617 => "010000110100001101000011",
14618 => "010000110100001101000011",
14619 => "010000110100001101000011",
14620 => "010000110100001101000011",
14621 => "010000110100001101000011",
14622 => "010011110100111101001111",
14623 => "011001100110011001100110",
14624 => "011001100110011001100110",
14625 => "010000110100001101000011",
14626 => "010000110100001101000011",
14627 => "010110100101101001011010",
14628 => "011001100110011001100110",
14629 => "010110110101101101011011",
14630 => "010000110100001101000011",
14631 => "010000110100001101000011",
14632 => "010000110100001101000011",
14633 => "010000110100001101000011",
14634 => "010000110100001101000011",
14635 => "010000110100001101000011",
14636 => "010000110100001101000011",
14637 => "010000110100001101000011",
14638 => "010000110100001101000011",
14639 => "011001100110011001100110",
14640 => "011001100110011001100110",
14641 => "010100010101000101010001",
14642 => "010000110100001101000011",
14643 => "010000110100001101000011",
14644 => "010000110100001101000011",
14645 => "010000110100001101000011",
14646 => "011001010110010101100101",
14647 => "011001100110011001100110",
14648 => "010100100101001001010010",
14649 => "010000110100001101000011",
14650 => "010000110100001101000011",
14651 => "010000110100001101000011",
14652 => "010000110100001101000011",
14653 => "010000110100001101000011",
14654 => "010000110100001101000011",
14655 => "010000110100001101000011",
14656 => "010000110100001101000011",
14657 => "010000110100001101000011",
14658 => "010000110100001101000011",
14659 => "010000110100001101000011",
14660 => "010000110100001101000011",
14661 => "010000110100001101000011",
14662 => "010000110100001101000011",
14663 => "010000110100001101000011",
14664 => "010000110100001101000011",
14665 => "010000110100001101000011",
14666 => "010000110100001101000011",
14667 => "010000110100001101000011",
14668 => "010000110100001101000011",
14669 => "010000110100001101000011",
14670 => "010000110100001101000011",
14671 => "001110110011101100111011",
14672 => "000000000000000000000000",
14673 => "000000000000000000000000",
14674 => "000000000000000000000000",
14675 => "000000000000000000000000",
14676 => "000000000000000000000000",
14677 => "000000000000000000000000",
14678 => "000000000000000000000000",
14679 => "000000000000000000000000",
14680 => "000000000000000000000000",
14681 => "000000000000000000000000",
14682 => "000000000000000000000000",
14683 => "000000000000000000000000",
14684 => "000000000000000000000000",
14685 => "000000000000000000000000",
14686 => "000000000000000000000000",
14687 => "000000000000000000000000",
14688 => "000000000000000000000000",
14689 => "000000000000000000000000",
14690 => "000000000000000000000000",
14691 => "000000000000000000000000",
14692 => "000000000000000000000000",
14693 => "000000000000000000000000",
14694 => "000000000000000000000000",
14695 => "000000000000000000000000",
14696 => "000000000000000000000000",
14697 => "000000000000000000000000",
14698 => "000000000000000000000000",
14699 => "000000000000000000000000",
14700 => "000000000000000000000000",
14701 => "000000000000000000000000",
14702 => "000000000000000000000000",
14703 => "000000000000000000000000",
14704 => "000000000000000000000000",
14705 => "000000000000000000000000",
14706 => "000000000000000000000000",
14707 => "000000000000000000000000",
14708 => "000000000000000000000000",
14709 => "000000000000000000000000",
14710 => "000000000000000000000000",
14711 => "000010110000101100001011",
14712 => "001001100010011000100110",
14713 => "001001100010011000100110",
14714 => "001001100010011000100110",
14715 => "001001100010011000100110",
14716 => "001101110011011100110111",
14717 => "010000110100001101000011",
14718 => "010000110100001101000011",
14719 => "010000110100001101000011",
14720 => "010000110100001101000011",
14721 => "010000110100001101000011",
14722 => "010000110100001101000011",
14723 => "010000110100001101000011",
14724 => "010000110100001101000011",
14725 => "010000110100001101000011",
14726 => "010000110100001101000011",
14727 => "010000110100001101000011",
14728 => "010000110100001101000011",
14729 => "010000110100001101000011",
14730 => "010000110100001101000011",
14731 => "010000110100001101000011",
14732 => "010000110100001101000011",
14733 => "010000110100001101000011",
14734 => "010000110100001101000011",
14735 => "010000110100001101000011",
14736 => "010000110100001101000011",
14737 => "010000110100001101000011",
14738 => "010000110100001101000011",
14739 => "010001010100010101000101",
14740 => "010100100101001001010010",
14741 => "010100100101001001010010",
14742 => "010001010100010101000101",
14743 => "010000110100001101000011",
14744 => "010000110100001101000011",
14745 => "010000110100001101000011",
14746 => "010001010100010101000101",
14747 => "010100100101001001010010",
14748 => "010100100101001001010010",
14749 => "010001100100011001000110",
14750 => "010000110100001101000011",
14751 => "010000110100001101000011",
14752 => "010000110100001101000011",
14753 => "010000110100001101000011",
14754 => "010000110100001101000011",
14755 => "010000110100001101000011",
14756 => "010100100101001001010010",
14757 => "010101110101011101010111",
14758 => "010101010101010101010101",
14759 => "010100100101001001010010",
14760 => "010100010101000101010001",
14761 => "010000110100001101000011",
14762 => "010000110100001101000011",
14763 => "010011100100111001001110",
14764 => "010100100101001001010010",
14765 => "010101000101010001010100",
14766 => "010101110101011101010111",
14767 => "010101100101011001010110",
14768 => "010000110100001101000011",
14769 => "010000110100001101000011",
14770 => "010100010101000101010001",
14771 => "010101110101011101010111",
14772 => "010101010101010101010101",
14773 => "010100100101001001010010",
14774 => "010100100101001001010010",
14775 => "010000110100001101000011",
14776 => "010000110100001101000011",
14777 => "010011010100110101001101",
14778 => "010100100101001001010010",
14779 => "010101000101010001010100",
14780 => "010101110101011101010111",
14781 => "010101110101011101010111",
14782 => "010000110100001101000011",
14783 => "010000110100001101000011",
14784 => "010000110100001101000011",
14785 => "010000110100001101000011",
14786 => "010000110100001101000011",
14787 => "010000110100001101000011",
14788 => "010000110100001101000011",
14789 => "010100100101001001010010",
14790 => "010100100101001001010010",
14791 => "010010010100100101001001",
14792 => "010000110100001101000011",
14793 => "010000110100001101000011",
14794 => "010000110100001101000011",
14795 => "010000110100001101000011",
14796 => "010100100101001001010010",
14797 => "010100100101001001010010",
14798 => "010010100100101001001010",
14799 => "010000110100001101000011",
14800 => "010000110100001101000011",
14801 => "010000110100001101000011",
14802 => "010000110100001101000011",
14803 => "010000110100001101000011",
14804 => "010000110100001101000011",
14805 => "010000110100001101000011",
14806 => "010000110100001101000011",
14807 => "010000110100001101000011",
14808 => "010000110100001101000011",
14809 => "010000110100001101000011",
14810 => "010000110100001101000011",
14811 => "010000110100001101000011",
14812 => "010000110100001101000011",
14813 => "010000110100001101000011",
14814 => "010000110100001101000011",
14815 => "010000110100001101000011",
14816 => "010000110100001101000011",
14817 => "010000110100001101000011",
14818 => "010000110100001101000011",
14819 => "010000110100001101000011",
14820 => "010000110100001101000011",
14821 => "001111110011111100111111",
14822 => "001001100010011000100110",
14823 => "001001100010011000100110",
14824 => "001001100010011000100110",
14825 => "001001100010011000100110",
14826 => "000101010001010100010101",
14827 => "000000000000000000000000",
14828 => "000000000000000000000000",
14829 => "000000000000000000000000",
14830 => "000000000000000000000000",
14831 => "000000000000000000000000",
14832 => "000000000000000000000000",
14833 => "000000000000000000000000",
14834 => "000000000000000000000000",
14835 => "000000000000000000000000",
14836 => "000000000000000000000000",
14837 => "000000000000000000000000",
14838 => "000000000000000000000000",
14839 => "000000000000000000000000",
14840 => "000000000000000000000000",
14841 => "000000000000000000000000",
14842 => "000000000000000000000000",
14843 => "000000000000000000000000",
14844 => "000000000000000000000000",
14845 => "000000000000000000000000",
14846 => "000000000000000000000000",
14847 => "000000000000000000000000",
14848 => "000000000000000000000000",
14849 => "000000000000000000000000",
14850 => "000000000000000000000000",
14851 => "000000000000000000000000",
14852 => "000000000000000000000000",
14853 => "000000000000000000000000",
14854 => "000000000000000000000000",
14855 => "000000000000000000000000",
14856 => "000000000000000000000000",
14857 => "000000000000000000000000",
14858 => "000000000000000000000000",
14859 => "000000000000000000000000",
14860 => "000000000000000000000000",
14861 => "000100110001001100010011",
14862 => "010000110100001101000011",
14863 => "010000110100001101000011",
14864 => "010000110100001101000011",
14865 => "010000110100001101000011",
14866 => "010000110100001101000011",
14867 => "010000110100001101000011",
14868 => "010000110100001101000011",
14869 => "010000110100001101000011",
14870 => "010000110100001101000011",
14871 => "010000110100001101000011",
14872 => "010000110100001101000011",
14873 => "010000110100001101000011",
14874 => "010000110100001101000011",
14875 => "010000110100001101000011",
14876 => "010000110100001101000011",
14877 => "010000110100001101000011",
14878 => "010000110100001101000011",
14879 => "010000110100001101000011",
14880 => "010000110100001101000011",
14881 => "010000110100001101000011",
14882 => "010000110100001101000011",
14883 => "010000110100001101000011",
14884 => "010000110100001101000011",
14885 => "010000110100001101000011",
14886 => "010000110100001101000011",
14887 => "010000110100001101000011",
14888 => "010000110100001101000011",
14889 => "010000110100001101000011",
14890 => "010000110100001101000011",
14891 => "010000110100001101000011",
14892 => "010000110100001101000011",
14893 => "010000110100001101000011",
14894 => "010000110100001101000011",
14895 => "010000110100001101000011",
14896 => "010000110100001101000011",
14897 => "010000110100001101000011",
14898 => "010000110100001101000011",
14899 => "010000110100001101000011",
14900 => "010000110100001101000011",
14901 => "010000110100001101000011",
14902 => "010000110100001101000011",
14903 => "010000110100001101000011",
14904 => "010000110100001101000011",
14905 => "010000110100001101000011",
14906 => "010111110101111101011111",
14907 => "011001100110011001100110",
14908 => "010110000101100001011000",
14909 => "010000110100001101000011",
14910 => "010000110100001101000011",
14911 => "010000110100001101000011",
14912 => "010000110100001101000011",
14913 => "010000110100001101000011",
14914 => "010000110100001101000011",
14915 => "010100000101000001010000",
14916 => "011001100110011001100110",
14917 => "011001010110010101100101",
14918 => "010000110100001101000011",
14919 => "010000110100001101000011",
14920 => "010110110101101101011011",
14921 => "011001100110011001100110",
14922 => "010110100101101001011010",
14923 => "010000110100001101000011",
14924 => "010000110100001101000011",
14925 => "010000110100001101000011",
14926 => "010000110100001101000011",
14927 => "010000110100001101000011",
14928 => "010000110100001101000011",
14929 => "010011100100111001001110",
14930 => "011001100110011001100110",
14931 => "011001100110011001100110",
14932 => "010000110100001101000011",
14933 => "010000110100001101000011",
14934 => "010000110100001101000011",
14935 => "010000110100001101000011",
14936 => "010000110100001101000011",
14937 => "010000110100001101000011",
14938 => "010000110100001101000011",
14939 => "010000110100001101000011",
14940 => "010000110100001101000011",
14941 => "010000110100001101000011",
14942 => "010000110100001101000011",
14943 => "010000110100001101000011",
14944 => "010000110100001101000011",
14945 => "010000110100001101000011",
14946 => "010000110100001101000011",
14947 => "010000110100001101000011",
14948 => "010000110100001101000011",
14949 => "010000110100001101000011",
14950 => "010000110100001101000011",
14951 => "010000110100001101000011",
14952 => "010000110100001101000011",
14953 => "010000110100001101000011",
14954 => "010000110100001101000011",
14955 => "010000110100001101000011",
14956 => "010000110100001101000011",
14957 => "010000110100001101000011",
14958 => "010000110100001101000011",
14959 => "010000110100001101000011",
14960 => "010000110100001101000011",
14961 => "010000110100001101000011",
14962 => "010000110100001101000011",
14963 => "010000110100001101000011",
14964 => "010000110100001101000011",
14965 => "010000110100001101000011",
14966 => "010000110100001101000011",
14967 => "010000110100001101000011",
14968 => "010000110100001101000011",
14969 => "010000110100001101000011",
14970 => "010000110100001101000011",
14971 => "010000110100001101000011",
14972 => "010000110100001101000011",
14973 => "010000110100001101000011",
14974 => "010000110100001101000011",
14975 => "010000110100001101000011",
14976 => "001001100010011000100110",
14977 => "000000000000000000000000",
14978 => "000000000000000000000000",
14979 => "000000000000000000000000",
14980 => "000000000000000000000000",
14981 => "000000000000000000000000",
14982 => "000000000000000000000000",
14983 => "000000000000000000000000",
14984 => "000000000000000000000000",
14985 => "000000000000000000000000",
14986 => "000000000000000000000000",
14987 => "000000000000000000000000",
14988 => "000000000000000000000000",
14989 => "000000000000000000000000",
14990 => "000000000000000000000000",
14991 => "000000000000000000000000",
14992 => "000000000000000000000000",
14993 => "000000000000000000000000",
14994 => "000000000000000000000000",
14995 => "000000000000000000000000",
14996 => "000000000000000000000000",
14997 => "000000000000000000000000",
14998 => "000000000000000000000000",
14999 => "000000000000000000000000",
15000 => "000000000000000000000000",
15001 => "000000000000000000000000",
15002 => "000000000000000000000000",
15003 => "000000000000000000000000",
15004 => "000000000000000000000000",
15005 => "000000000000000000000000",
15006 => "000000000000000000000000",
15007 => "000000000000000000000000",
15008 => "000000000000000000000000",
15009 => "000000000000000000000000",
15010 => "000000000000000000000000",
15011 => "000100110001001100010011",
15012 => "010000110100001101000011",
15013 => "010000110100001101000011",
15014 => "010000110100001101000011",
15015 => "010000110100001101000011",
15016 => "010000110100001101000011",
15017 => "010000110100001101000011",
15018 => "010000110100001101000011",
15019 => "010000110100001101000011",
15020 => "010000110100001101000011",
15021 => "010000110100001101000011",
15022 => "010000110100001101000011",
15023 => "010000110100001101000011",
15024 => "010000110100001101000011",
15025 => "010000110100001101000011",
15026 => "010000110100001101000011",
15027 => "010000110100001101000011",
15028 => "010000110100001101000011",
15029 => "010000110100001101000011",
15030 => "010000110100001101000011",
15031 => "010000110100001101000011",
15032 => "010000110100001101000011",
15033 => "010000110100001101000011",
15034 => "010000110100001101000011",
15035 => "010000110100001101000011",
15036 => "010000110100001101000011",
15037 => "010000110100001101000011",
15038 => "010000110100001101000011",
15039 => "010000110100001101000011",
15040 => "010000110100001101000011",
15041 => "010000110100001101000011",
15042 => "010000110100001101000011",
15043 => "010000110100001101000011",
15044 => "010000110100001101000011",
15045 => "010000110100001101000011",
15046 => "010000110100001101000011",
15047 => "010000110100001101000011",
15048 => "010000110100001101000011",
15049 => "010000110100001101000011",
15050 => "010000110100001101000011",
15051 => "010000110100001101000011",
15052 => "010000110100001101000011",
15053 => "010000110100001101000011",
15054 => "010000110100001101000011",
15055 => "010000110100001101000011",
15056 => "010111110101111101011111",
15057 => "011001100110011001100110",
15058 => "010110000101100001011000",
15059 => "010000110100001101000011",
15060 => "010000110100001101000011",
15061 => "010000110100001101000011",
15062 => "010000110100001101000011",
15063 => "010000110100001101000011",
15064 => "010000110100001101000011",
15065 => "010100000101000001010000",
15066 => "011001100110011001100110",
15067 => "011001010110010101100101",
15068 => "010000110100001101000011",
15069 => "010000110100001101000011",
15070 => "010110110101101101011011",
15071 => "011001100110011001100110",
15072 => "010110100101101001011010",
15073 => "010000110100001101000011",
15074 => "010000110100001101000011",
15075 => "010000110100001101000011",
15076 => "010000110100001101000011",
15077 => "010000110100001101000011",
15078 => "010000110100001101000011",
15079 => "010011100100111001001110",
15080 => "011001100110011001100110",
15081 => "011001100110011001100110",
15082 => "010000110100001101000011",
15083 => "010000110100001101000011",
15084 => "010000110100001101000011",
15085 => "010000110100001101000011",
15086 => "010000110100001101000011",
15087 => "010000110100001101000011",
15088 => "010000110100001101000011",
15089 => "010000110100001101000011",
15090 => "010000110100001101000011",
15091 => "010000110100001101000011",
15092 => "010000110100001101000011",
15093 => "010000110100001101000011",
15094 => "010000110100001101000011",
15095 => "010000110100001101000011",
15096 => "010000110100001101000011",
15097 => "010000110100001101000011",
15098 => "010000110100001101000011",
15099 => "010000110100001101000011",
15100 => "010000110100001101000011",
15101 => "010000110100001101000011",
15102 => "010000110100001101000011",
15103 => "010000110100001101000011",
15104 => "010000110100001101000011",
15105 => "010000110100001101000011",
15106 => "010000110100001101000011",
15107 => "010000110100001101000011",
15108 => "010000110100001101000011",
15109 => "010000110100001101000011",
15110 => "010000110100001101000011",
15111 => "010000110100001101000011",
15112 => "010000110100001101000011",
15113 => "010000110100001101000011",
15114 => "010000110100001101000011",
15115 => "010000110100001101000011",
15116 => "010000110100001101000011",
15117 => "010000110100001101000011",
15118 => "010000110100001101000011",
15119 => "010000110100001101000011",
15120 => "010000110100001101000011",
15121 => "010000110100001101000011",
15122 => "010000110100001101000011",
15123 => "010000110100001101000011",
15124 => "010000110100001101000011",
15125 => "010000110100001101000011",
15126 => "001001100010011000100110",
15127 => "000000000000000000000000",
15128 => "000000000000000000000000",
15129 => "000000000000000000000000",
15130 => "000000000000000000000000",
15131 => "000000000000000000000000",
15132 => "000000000000000000000000",
15133 => "000000000000000000000000",
15134 => "000000000000000000000000",
15135 => "000000000000000000000000",
15136 => "000000000000000000000000",
15137 => "000000000000000000000000",
15138 => "000000000000000000000000",
15139 => "000000000000000000000000",
15140 => "000000000000000000000000",
15141 => "000000000000000000000000",
15142 => "000000000000000000000000",
15143 => "000000000000000000000000",
15144 => "000000000000000000000000",
15145 => "000000000000000000000000",
15146 => "000000000000000000000000",
15147 => "000000000000000000000000",
15148 => "000000000000000000000000",
15149 => "000000000000000000000000",
15150 => "000000000000000000000000",
15151 => "000000000000000000000000",
15152 => "000000000000000000000000",
15153 => "000000000000000000000000",
15154 => "000000000000000000000000",
15155 => "000000000000000000000000",
15156 => "000000000000000000000000",
15157 => "000000000000000000000000",
15158 => "000000000000000000000000",
15159 => "000000000000000000000000",
15160 => "000000000000000000000000",
15161 => "000100110001001100010011",
15162 => "010000110100001101000011",
15163 => "010000110100001101000011",
15164 => "010000110100001101000011",
15165 => "010000110100001101000011",
15166 => "010000110100001101000011",
15167 => "010000110100001101000011",
15168 => "010000110100001101000011",
15169 => "010000110100001101000011",
15170 => "010000110100001101000011",
15171 => "010000110100001101000011",
15172 => "010000110100001101000011",
15173 => "010000110100001101000011",
15174 => "010000110100001101000011",
15175 => "010000110100001101000011",
15176 => "010000110100001101000011",
15177 => "010000110100001101000011",
15178 => "010000110100001101000011",
15179 => "010000110100001101000011",
15180 => "010000110100001101000011",
15181 => "010000110100001101000011",
15182 => "010000110100001101000011",
15183 => "010000110100001101000011",
15184 => "010000110100001101000011",
15185 => "010000110100001101000011",
15186 => "010000110100001101000011",
15187 => "010000110100001101000011",
15188 => "010000110100001101000011",
15189 => "010000110100001101000011",
15190 => "010000110100001101000011",
15191 => "010000110100001101000011",
15192 => "010000110100001101000011",
15193 => "010000110100001101000011",
15194 => "010000110100001101000011",
15195 => "010000110100001101000011",
15196 => "010000110100001101000011",
15197 => "010000110100001101000011",
15198 => "010000110100001101000011",
15199 => "010000110100001101000011",
15200 => "010000110100001101000011",
15201 => "010000110100001101000011",
15202 => "010000110100001101000011",
15203 => "010000110100001101000011",
15204 => "010000110100001101000011",
15205 => "010000110100001101000011",
15206 => "010111110101111101011111",
15207 => "011001100110011001100110",
15208 => "010110000101100001011000",
15209 => "010000110100001101000011",
15210 => "010000110100001101000011",
15211 => "010000110100001101000011",
15212 => "010000110100001101000011",
15213 => "010000110100001101000011",
15214 => "010000110100001101000011",
15215 => "010100000101000001010000",
15216 => "011001100110011001100110",
15217 => "011001010110010101100101",
15218 => "010000110100001101000011",
15219 => "010000110100001101000011",
15220 => "010110110101101101011011",
15221 => "011001100110011001100110",
15222 => "010110100101101001011010",
15223 => "010000110100001101000011",
15224 => "010000110100001101000011",
15225 => "010000110100001101000011",
15226 => "010000110100001101000011",
15227 => "010000110100001101000011",
15228 => "010000110100001101000011",
15229 => "010011100100111001001110",
15230 => "011001100110011001100110",
15231 => "011001100110011001100110",
15232 => "010000110100001101000011",
15233 => "010000110100001101000011",
15234 => "010000110100001101000011",
15235 => "010000110100001101000011",
15236 => "010000110100001101000011",
15237 => "010000110100001101000011",
15238 => "010000110100001101000011",
15239 => "010000110100001101000011",
15240 => "010000110100001101000011",
15241 => "010000110100001101000011",
15242 => "010000110100001101000011",
15243 => "010000110100001101000011",
15244 => "010000110100001101000011",
15245 => "010000110100001101000011",
15246 => "010000110100001101000011",
15247 => "010000110100001101000011",
15248 => "010000110100001101000011",
15249 => "010000110100001101000011",
15250 => "010000110100001101000011",
15251 => "010000110100001101000011",
15252 => "010000110100001101000011",
15253 => "010000110100001101000011",
15254 => "010000110100001101000011",
15255 => "010000110100001101000011",
15256 => "010000110100001101000011",
15257 => "010000110100001101000011",
15258 => "010000110100001101000011",
15259 => "010000110100001101000011",
15260 => "010000110100001101000011",
15261 => "010000110100001101000011",
15262 => "010000110100001101000011",
15263 => "010000110100001101000011",
15264 => "010000110100001101000011",
15265 => "010000110100001101000011",
15266 => "010000110100001101000011",
15267 => "010000110100001101000011",
15268 => "010000110100001101000011",
15269 => "010000110100001101000011",
15270 => "010000110100001101000011",
15271 => "010000110100001101000011",
15272 => "010000110100001101000011",
15273 => "010000110100001101000011",
15274 => "010000110100001101000011",
15275 => "010000110100001101000011",
15276 => "001001100010011000100110",
15277 => "000000000000000000000000",
15278 => "000000000000000000000000",
15279 => "000000000000000000000000",
15280 => "000000000000000000000000",
15281 => "000000000000000000000000",
15282 => "000000000000000000000000",
15283 => "000000000000000000000000",
15284 => "000000000000000000000000",
15285 => "000000000000000000000000",
15286 => "000000000000000000000000",
15287 => "000000000000000000000000",
15288 => "000000000000000000000000",
15289 => "000000000000000000000000",
15290 => "000000000000000000000000",
15291 => "000000000000000000000000",
15292 => "000000000000000000000000",
15293 => "000000000000000000000000",
15294 => "000000000000000000000000",
15295 => "000000000000000000000000",
15296 => "000000000000000000000000",
15297 => "000000000000000000000000",
15298 => "000000000000000000000000",
15299 => "000000000000000000000000",
15300 => "000000000000000000000000",
15301 => "000000000000000000000000",
15302 => "000000000000000000000000",
15303 => "000000000000000000000000",
15304 => "000000000000000000000000",
15305 => "000000000000000000000000",
15306 => "000000000000000000000000",
15307 => "000000000000000000000000",
15308 => "000000000000000000000000",
15309 => "000000000000000000000000",
15310 => "000000000000000000000000",
15311 => "000100110001001100010011",
15312 => "010000110100001101000011",
15313 => "010000110100001101000011",
15314 => "010000110100001101000011",
15315 => "010000110100001101000011",
15316 => "010000110100001101000011",
15317 => "010000110100001101000011",
15318 => "010000110100001101000011",
15319 => "010000110100001101000011",
15320 => "010000110100001101000011",
15321 => "010000110100001101000011",
15322 => "010000110100001101000011",
15323 => "010000110100001101000011",
15324 => "010000110100001101000011",
15325 => "010000110100001101000011",
15326 => "010000110100001101000011",
15327 => "010000110100001101000011",
15328 => "010000110100001101000011",
15329 => "010000110100001101000011",
15330 => "010000110100001101000011",
15331 => "010000110100001101000011",
15332 => "010000110100001101000011",
15333 => "010000110100001101000011",
15334 => "010000110100001101000011",
15335 => "010000110100001101000011",
15336 => "010000110100001101000011",
15337 => "010000110100001101000011",
15338 => "010000110100001101000011",
15339 => "010000110100001101000011",
15340 => "010000110100001101000011",
15341 => "010000110100001101000011",
15342 => "010000110100001101000011",
15343 => "010000110100001101000011",
15344 => "010000110100001101000011",
15345 => "010000110100001101000011",
15346 => "010000110100001101000011",
15347 => "010000110100001101000011",
15348 => "010000110100001101000011",
15349 => "010000110100001101000011",
15350 => "010000110100001101000011",
15351 => "010000110100001101000011",
15352 => "010000110100001101000011",
15353 => "010000110100001101000011",
15354 => "010000110100001101000011",
15355 => "010000110100001101000011",
15356 => "010111110101111101011111",
15357 => "011001100110011001100110",
15358 => "010110000101100001011000",
15359 => "010000110100001101000011",
15360 => "010000110100001101000011",
15361 => "010000110100001101000011",
15362 => "010000110100001101000011",
15363 => "010000110100001101000011",
15364 => "010000110100001101000011",
15365 => "010100000101000001010000",
15366 => "011001100110011001100110",
15367 => "011001010110010101100101",
15368 => "010000110100001101000011",
15369 => "010000110100001101000011",
15370 => "010110110101101101011011",
15371 => "011001100110011001100110",
15372 => "010110100101101001011010",
15373 => "010000110100001101000011",
15374 => "010000110100001101000011",
15375 => "010000110100001101000011",
15376 => "010000110100001101000011",
15377 => "010000110100001101000011",
15378 => "010000110100001101000011",
15379 => "010011100100111001001110",
15380 => "011001100110011001100110",
15381 => "011001100110011001100110",
15382 => "010000110100001101000011",
15383 => "010000110100001101000011",
15384 => "010000110100001101000011",
15385 => "010000110100001101000011",
15386 => "010000110100001101000011",
15387 => "010000110100001101000011",
15388 => "010000110100001101000011",
15389 => "010000110100001101000011",
15390 => "010000110100001101000011",
15391 => "010000110100001101000011",
15392 => "010000110100001101000011",
15393 => "010000110100001101000011",
15394 => "010000110100001101000011",
15395 => "010000110100001101000011",
15396 => "010000110100001101000011",
15397 => "010000110100001101000011",
15398 => "010000110100001101000011",
15399 => "010000110100001101000011",
15400 => "010000110100001101000011",
15401 => "010000110100001101000011",
15402 => "010000110100001101000011",
15403 => "010000110100001101000011",
15404 => "010000110100001101000011",
15405 => "010000110100001101000011",
15406 => "010000110100001101000011",
15407 => "010000110100001101000011",
15408 => "010000110100001101000011",
15409 => "010000110100001101000011",
15410 => "010000110100001101000011",
15411 => "010000110100001101000011",
15412 => "010000110100001101000011",
15413 => "010000110100001101000011",
15414 => "010000110100001101000011",
15415 => "010000110100001101000011",
15416 => "010000110100001101000011",
15417 => "010000110100001101000011",
15418 => "010000110100001101000011",
15419 => "010000110100001101000011",
15420 => "010000110100001101000011",
15421 => "010000110100001101000011",
15422 => "010000110100001101000011",
15423 => "010000110100001101000011",
15424 => "010000110100001101000011",
15425 => "010000110100001101000011",
15426 => "001001100010011000100110",
15427 => "000000000000000000000000",
15428 => "000000000000000000000000",
15429 => "000000000000000000000000",
15430 => "000000000000000000000000",
15431 => "000000000000000000000000",
15432 => "000000000000000000000000",
15433 => "000000000000000000000000",
15434 => "000000000000000000000000",
15435 => "000000000000000000000000",
15436 => "000000000000000000000000",
15437 => "000000000000000000000000",
15438 => "000000000000000000000000",
15439 => "000000000000000000000000",
15440 => "000000000000000000000000",
15441 => "000000000000000000000000",
15442 => "000000000000000000000000",
15443 => "000000000000000000000000",
15444 => "000000000000000000000000",
15445 => "000000000000000000000000",
15446 => "000000000000000000000000",
15447 => "000000000000000000000000",
15448 => "000000000000000000000000",
15449 => "000000000000000000000000",
15450 => "000000000000000000000000",
15451 => "000000000000000000000000",
15452 => "000000000000000000000000",
15453 => "000000000000000000000000",
15454 => "000000000000000000000000",
15455 => "000000000000000000000000",
15456 => "000000000000000000000000",
15457 => "000000000000000000000000",
15458 => "000000000000000000000000",
15459 => "000000000000000000000000",
15460 => "000000000000000000000000",
15461 => "000000010000000100000001",
15462 => "000001000000010000000100",
15463 => "000001000000010000000100",
15464 => "010000100100001001000010",
15465 => "010000110100001101000011",
15466 => "010000110100001101000011",
15467 => "010000110100001101000011",
15468 => "010000110100001101000011",
15469 => "010000110100001101000011",
15470 => "010000110100001101000011",
15471 => "010000110100001101000011",
15472 => "010000110100001101000011",
15473 => "010000110100001101000011",
15474 => "010000110100001101000011",
15475 => "010000110100001101000011",
15476 => "010000110100001101000011",
15477 => "010000110100001101000011",
15478 => "010000110100001101000011",
15479 => "010000110100001101000011",
15480 => "001000010010000100100001",
15481 => "000001000000010000000100",
15482 => "000001000000010000000100",
15483 => "000001000000010000000100",
15484 => "000001000000010000000100",
15485 => "000001000000010000000100",
15486 => "000001000000010000000100",
15487 => "000001000000010000000100",
15488 => "000001000000010000000100",
15489 => "000001000000010000000100",
15490 => "000001000000010000000100",
15491 => "000001000000010000000100",
15492 => "000001000000010000000100",
15493 => "000001000000010000000100",
15494 => "000001000000010000000100",
15495 => "000001000000010000000100",
15496 => "000001000000010000000100",
15497 => "000001000000010000000100",
15498 => "000001000000010000000100",
15499 => "000001000000010000000100",
15500 => "000001000000010000000100",
15501 => "000001000000010000000100",
15502 => "000001000000010000000100",
15503 => "000010100000101000001010",
15504 => "010000110100001101000011",
15505 => "010000110100001101000011",
15506 => "010111110101111101011111",
15507 => "011001100110011001100110",
15508 => "010110000101100001011000",
15509 => "010000110100001101000011",
15510 => "010000110100001101000011",
15511 => "010000110100001101000011",
15512 => "010000110100001101000011",
15513 => "010000110100001101000011",
15514 => "010000110100001101000011",
15515 => "010100000101000001010000",
15516 => "011001100110011001100110",
15517 => "011001010110010101100101",
15518 => "010000110100001101000011",
15519 => "010000110100001101000011",
15520 => "010110110101101101011011",
15521 => "011001100110011001100110",
15522 => "010110100101101001011010",
15523 => "010000110100001101000011",
15524 => "010000110100001101000011",
15525 => "010000110100001101000011",
15526 => "010000110100001101000011",
15527 => "010000110100001101000011",
15528 => "010000110100001101000011",
15529 => "010011100100111001001110",
15530 => "011001100110011001100110",
15531 => "011001100110011001100110",
15532 => "010000110100001101000011",
15533 => "010000110100001101000011",
15534 => "000110110001101100011011",
15535 => "000001000000010000000100",
15536 => "000001000000010000000100",
15537 => "000001000000010000000100",
15538 => "000001000000010000000100",
15539 => "000001000000010000000100",
15540 => "000001000000010000000100",
15541 => "000001000000010000000100",
15542 => "000001000000010000000100",
15543 => "000001000000010000000100",
15544 => "000001000000010000000100",
15545 => "000001000000010000000100",
15546 => "000001000000010000000100",
15547 => "000001000000010000000100",
15548 => "000001000000010000000100",
15549 => "000001000000010000000100",
15550 => "000001000000010000000100",
15551 => "000001000000010000000100",
15552 => "000001000000010000000100",
15553 => "000001000000010000000100",
15554 => "000001000000010000000100",
15555 => "000001000000010000000100",
15556 => "000001000000010000000100",
15557 => "000011110000111100001111",
15558 => "010000110100001101000011",
15559 => "010000110100001101000011",
15560 => "010000110100001101000011",
15561 => "010000110100001101000011",
15562 => "010000110100001101000011",
15563 => "010000110100001101000011",
15564 => "010000110100001101000011",
15565 => "010000110100001101000011",
15566 => "010000110100001101000011",
15567 => "010000110100001101000011",
15568 => "010000110100001101000011",
15569 => "010000110100001101000011",
15570 => "010000110100001101000011",
15571 => "010000110100001101000011",
15572 => "010000110100001101000011",
15573 => "010000110100001101000011",
15574 => "000011100000111000001110",
15575 => "000001000000010000000100",
15576 => "000000100000001000000010",
15577 => "000000000000000000000000",
15578 => "000000000000000000000000",
15579 => "000000000000000000000000",
15580 => "000000000000000000000000",
15581 => "000000000000000000000000",
15582 => "000000000000000000000000",
15583 => "000000000000000000000000",
15584 => "000000000000000000000000",
15585 => "000000000000000000000000",
15586 => "000000000000000000000000",
15587 => "000000000000000000000000",
15588 => "000000000000000000000000",
15589 => "000000000000000000000000",
15590 => "000000000000000000000000",
15591 => "000000000000000000000000",
15592 => "000000000000000000000000",
15593 => "000000000000000000000000",
15594 => "000000000000000000000000",
15595 => "000000000000000000000000",
15596 => "000000000000000000000000",
15597 => "000000000000000000000000",
15598 => "000000000000000000000000",
15599 => "000000000000000000000000",
15600 => "000000000000000000000000",
15601 => "000000000000000000000000",
15602 => "000000000000000000000000",
15603 => "000000000000000000000000",
15604 => "000000000000000000000000",
15605 => "000000000000000000000000",
15606 => "000000000000000000000000",
15607 => "000000000000000000000000",
15608 => "000000000000000000000000",
15609 => "000000000000000000000000",
15610 => "000000000000000000000000",
15611 => "000000000000000000000000",
15612 => "000000000000000000000000",
15613 => "000000000000000000000000",
15614 => "010000100100001001000010",
15615 => "010000110100001101000011",
15616 => "010000110100001101000011",
15617 => "010000110100001101000011",
15618 => "010000110100001101000011",
15619 => "010000110100001101000011",
15620 => "010000110100001101000011",
15621 => "010000110100001101000011",
15622 => "010000110100001101000011",
15623 => "010000110100001101000011",
15624 => "010000110100001101000011",
15625 => "010000110100001101000011",
15626 => "010000110100001101000011",
15627 => "010000110100001101000011",
15628 => "010000110100001101000011",
15629 => "010000110100001101000011",
15630 => "000111110001111100011111",
15631 => "000000000000000000000000",
15632 => "000000000000000000000000",
15633 => "000000000000000000000000",
15634 => "000000000000000000000000",
15635 => "000000000000000000000000",
15636 => "000000000000000000000000",
15637 => "000000000000000000000000",
15638 => "000000000000000000000000",
15639 => "000000000000000000000000",
15640 => "000000000000000000000000",
15641 => "000000000000000000000000",
15642 => "000000000000000000000000",
15643 => "000000000000000000000000",
15644 => "000000000000000000000000",
15645 => "000000000000000000000000",
15646 => "000000000000000000000000",
15647 => "000000000000000000000000",
15648 => "000000000000000000000000",
15649 => "000000000000000000000000",
15650 => "000000000000000000000000",
15651 => "000000000000000000000000",
15652 => "000000000000000000000000",
15653 => "000001100000011000000110",
15654 => "010000110100001101000011",
15655 => "010000110100001101000011",
15656 => "010111110101111101011111",
15657 => "011001100110011001100110",
15658 => "010110000101100001011000",
15659 => "010000110100001101000011",
15660 => "010000110100001101000011",
15661 => "010000110100001101000011",
15662 => "010000110100001101000011",
15663 => "010000110100001101000011",
15664 => "010000110100001101000011",
15665 => "010100000101000001010000",
15666 => "011001100110011001100110",
15667 => "011001010110010101100101",
15668 => "010000110100001101000011",
15669 => "010000110100001101000011",
15670 => "010110110101101101011011",
15671 => "011001100110011001100110",
15672 => "010110100101101001011010",
15673 => "010000110100001101000011",
15674 => "010000110100001101000011",
15675 => "010000110100001101000011",
15676 => "010000110100001101000011",
15677 => "010000110100001101000011",
15678 => "010000110100001101000011",
15679 => "010011100100111001001110",
15680 => "011001100110011001100110",
15681 => "011001100110011001100110",
15682 => "010000110100001101000011",
15683 => "010000110100001101000011",
15684 => "000110010001100100011001",
15685 => "000000000000000000000000",
15686 => "000000000000000000000000",
15687 => "000000000000000000000000",
15688 => "000000000000000000000000",
15689 => "000000000000000000000000",
15690 => "000000000000000000000000",
15691 => "000000000000000000000000",
15692 => "000000000000000000000000",
15693 => "000000000000000000000000",
15694 => "000000000000000000000000",
15695 => "000000000000000000000000",
15696 => "000000000000000000000000",
15697 => "000000000000000000000000",
15698 => "000000000000000000000000",
15699 => "000000000000000000000000",
15700 => "000000000000000000000000",
15701 => "000000000000000000000000",
15702 => "000000000000000000000000",
15703 => "000000000000000000000000",
15704 => "000000000000000000000000",
15705 => "000000000000000000000000",
15706 => "000000000000000000000000",
15707 => "000011010000110100001101",
15708 => "010000110100001101000011",
15709 => "010000110100001101000011",
15710 => "010000110100001101000011",
15711 => "010000110100001101000011",
15712 => "010000110100001101000011",
15713 => "010000110100001101000011",
15714 => "010000110100001101000011",
15715 => "010000110100001101000011",
15716 => "010000110100001101000011",
15717 => "010000110100001101000011",
15718 => "010000110100001101000011",
15719 => "010000110100001101000011",
15720 => "010000110100001101000011",
15721 => "010000110100001101000011",
15722 => "010000110100001101000011",
15723 => "010000110100001101000011",
15724 => "000010110000101100001011",
15725 => "000000000000000000000000",
15726 => "000000000000000000000000",
15727 => "000000000000000000000000",
15728 => "000000000000000000000000",
15729 => "000000000000000000000000",
15730 => "000000000000000000000000",
15731 => "000000000000000000000000",
15732 => "000000000000000000000000",
15733 => "000000000000000000000000",
15734 => "000000000000000000000000",
15735 => "000000000000000000000000",
15736 => "000000000000000000000000",
15737 => "000000000000000000000000",
15738 => "000000000000000000000000",
15739 => "000000000000000000000000",
15740 => "000000000000000000000000",
15741 => "000000000000000000000000",
15742 => "000000000000000000000000",
15743 => "000000000000000000000000",
15744 => "000000000000000000000000",
15745 => "000000000000000000000000",
15746 => "000000000000000000000000",
15747 => "000000000000000000000000",
15748 => "000000000000000000000000",
15749 => "000000000000000000000000",
15750 => "000000000000000000000000",
15751 => "000000000000000000000000",
15752 => "000000000000000000000000",
15753 => "000000000000000000000000",
15754 => "000000000000000000000000",
15755 => "000000000000000000000000",
15756 => "000000000000000000000000",
15757 => "000000000000000000000000",
15758 => "000000000000000000000000",
15759 => "000000000000000000000000",
15760 => "000000000000000000000000",
15761 => "000000000000000000000000",
15762 => "000000000000000000000000",
15763 => "000000000000000000000000",
15764 => "010000100100001001000010",
15765 => "010000110100001101000011",
15766 => "010000110100001101000011",
15767 => "010000110100001101000011",
15768 => "001110100011101000111010",
15769 => "000111110001111100011111",
15770 => "000111110001111100011111",
15771 => "000111110001111100011111",
15772 => "000111110001111100011111",
15773 => "000111110001111100011111",
15774 => "000111110001111100011111",
15775 => "000111110001111100011111",
15776 => "000111110001111100011111",
15777 => "000111110001111100011111",
15778 => "000111110001111100011111",
15779 => "000111110001111100011111",
15780 => "000011110000111100001111",
15781 => "000000000000000000000000",
15782 => "000000000000000000000000",
15783 => "000000000000000000000000",
15784 => "000000000000000000000000",
15785 => "000000000000000000000000",
15786 => "000000000000000000000000",
15787 => "000000000000000000000000",
15788 => "000000000000000000000000",
15789 => "000000000000000000000000",
15790 => "000000000000000000000000",
15791 => "000000000000000000000000",
15792 => "000000000000000000000000",
15793 => "000000000000000000000000",
15794 => "000000000000000000000000",
15795 => "000000000000000000000000",
15796 => "000000000000000000000000",
15797 => "000000000000000000000000",
15798 => "000000000000000000000000",
15799 => "000000000000000000000000",
15800 => "000000000000000000000000",
15801 => "000000000000000000000000",
15802 => "000000000000000000000000",
15803 => "000000110000001100000011",
15804 => "000111110001111100011111",
15805 => "000111110001111100011111",
15806 => "010101110101011101010111",
15807 => "011001100110011001100110",
15808 => "010110000101100001011000",
15809 => "010000110100001101000011",
15810 => "010000110100001101000011",
15811 => "010000110100001101000011",
15812 => "010000110100001101000011",
15813 => "010000110100001101000011",
15814 => "010000110100001101000011",
15815 => "010100000101000001010000",
15816 => "011001100110011001100110",
15817 => "011001010110010101100101",
15818 => "010000110100001101000011",
15819 => "010000110100001101000011",
15820 => "010110110101101101011011",
15821 => "011001100110011001100110",
15822 => "010110100101101001011010",
15823 => "010000110100001101000011",
15824 => "010000110100001101000011",
15825 => "010000110100001101000011",
15826 => "010000110100001101000011",
15827 => "010000110100001101000011",
15828 => "010000110100001101000011",
15829 => "010011100100111001001110",
15830 => "011001100110011001100110",
15831 => "011001100110011001100110",
15832 => "001000000010000000100000",
15833 => "000111110001111100011111",
15834 => "000011000000110000001100",
15835 => "000000000000000000000000",
15836 => "000000000000000000000000",
15837 => "000000000000000000000000",
15838 => "000000000000000000000000",
15839 => "000000000000000000000000",
15840 => "000000000000000000000000",
15841 => "000000000000000000000000",
15842 => "000000000000000000000000",
15843 => "000000000000000000000000",
15844 => "000000000000000000000000",
15845 => "000000000000000000000000",
15846 => "000000000000000000000000",
15847 => "000000000000000000000000",
15848 => "000000000000000000000000",
15849 => "000000000000000000000000",
15850 => "000000000000000000000000",
15851 => "000000000000000000000000",
15852 => "000000000000000000000000",
15853 => "000000000000000000000000",
15854 => "000000000000000000000000",
15855 => "000000000000000000000000",
15856 => "000000000000000000000000",
15857 => "000001100000011000000110",
15858 => "000111110001111100011111",
15859 => "000111110001111100011111",
15860 => "000111110001111100011111",
15861 => "000111110001111100011111",
15862 => "000111110001111100011111",
15863 => "000111110001111100011111",
15864 => "000111110001111100011111",
15865 => "000111110001111100011111",
15866 => "000111110001111100011111",
15867 => "000111110001111100011111",
15868 => "000111110001111100011111",
15869 => "001100000011000000110000",
15870 => "010000110100001101000011",
15871 => "010000110100001101000011",
15872 => "010000110100001101000011",
15873 => "010000110100001101000011",
15874 => "000010110000101100001011",
15875 => "000000000000000000000000",
15876 => "000000000000000000000000",
15877 => "000000000000000000000000",
15878 => "000000000000000000000000",
15879 => "000000000000000000000000",
15880 => "000000000000000000000000",
15881 => "000000000000000000000000",
15882 => "000000000000000000000000",
15883 => "000000000000000000000000",
15884 => "000000000000000000000000",
15885 => "000000000000000000000000",
15886 => "000000000000000000000000",
15887 => "000000000000000000000000",
15888 => "000000000000000000000000",
15889 => "000000000000000000000000",
15890 => "000000000000000000000000",
15891 => "000000000000000000000000",
15892 => "000000000000000000000000",
15893 => "000000000000000000000000",
15894 => "000000000000000000000000",
15895 => "000000000000000000000000",
15896 => "000000000000000000000000",
15897 => "000000000000000000000000",
15898 => "000000000000000000000000",
15899 => "000000000000000000000000",
15900 => "000000000000000000000000",
15901 => "000000000000000000000000",
15902 => "000000000000000000000000",
15903 => "000000000000000000000000",
15904 => "000000000000000000000000",
15905 => "000000000000000000000000",
15906 => "000000000000000000000000",
15907 => "000000000000000000000000",
15908 => "000000000000000000000000",
15909 => "000000000000000000000000",
15910 => "000000000000000000000000",
15911 => "000000000000000000000000",
15912 => "000000000000000000000000",
15913 => "000000000000000000000000",
15914 => "010000100100001001000010",
15915 => "010000110100001101000011",
15916 => "010000110100001101000011",
15917 => "010000110100001101000011",
15918 => "001100100011001000110010",
15919 => "000000000000000000000000",
15920 => "000000000000000000000000",
15921 => "000000000000000000000000",
15922 => "000000000000000000000000",
15923 => "000000000000000000000000",
15924 => "000000000000000000000000",
15925 => "000000000000000000000000",
15926 => "000000000000000000000000",
15927 => "000000000000000000000000",
15928 => "000000000000000000000000",
15929 => "000000000000000000000000",
15930 => "000000000000000000000000",
15931 => "000000000000000000000000",
15932 => "000000000000000000000000",
15933 => "000000000000000000000000",
15934 => "000000000000000000000000",
15935 => "000000000000000000000000",
15936 => "000000000000000000000000",
15937 => "000000000000000000000000",
15938 => "000000000000000000000000",
15939 => "000000000000000000000000",
15940 => "000000000000000000000000",
15941 => "000000000000000000000000",
15942 => "000000000000000000000000",
15943 => "000000000000000000000000",
15944 => "000000000000000000000000",
15945 => "000000000000000000000000",
15946 => "000000000000000000000000",
15947 => "000000000000000000000000",
15948 => "000000000000000000000000",
15949 => "000000000000000000000000",
15950 => "000000000000000000000000",
15951 => "000000000000000000000000",
15952 => "000000000000000000000000",
15953 => "000000000000000000000000",
15954 => "000000000000000000000000",
15955 => "000000000000000000000000",
15956 => "010100000101000001010000",
15957 => "011001100110011001100110",
15958 => "010110000101100001011000",
15959 => "010000110100001101000011",
15960 => "010000110100001101000011",
15961 => "010000110100001101000011",
15962 => "010000110100001101000011",
15963 => "010000110100001101000011",
15964 => "010000110100001101000011",
15965 => "010100000101000001010000",
15966 => "011001100110011001100110",
15967 => "011001010110010101100101",
15968 => "010000110100001101000011",
15969 => "010000110100001101000011",
15970 => "010110110101101101011011",
15971 => "011001100110011001100110",
15972 => "010110100101101001011010",
15973 => "010000110100001101000011",
15974 => "010000110100001101000011",
15975 => "010000110100001101000011",
15976 => "010000110100001101000011",
15977 => "010000110100001101000011",
15978 => "010000110100001101000011",
15979 => "010011100100111001001110",
15980 => "011001100110011001100110",
15981 => "011001100110011001100110",
15982 => "000000000000000000000000",
15983 => "000000000000000000000000",
15984 => "000000000000000000000000",
15985 => "000000000000000000000000",
15986 => "000000000000000000000000",
15987 => "000000000000000000000000",
15988 => "000000000000000000000000",
15989 => "000000000000000000000000",
15990 => "000000000000000000000000",
15991 => "000000000000000000000000",
15992 => "000000000000000000000000",
15993 => "000000000000000000000000",
15994 => "000000000000000000000000",
15995 => "000000000000000000000000",
15996 => "000000000000000000000000",
15997 => "000000000000000000000000",
15998 => "000000000000000000000000",
15999 => "000000000000000000000000",
16000 => "000000000000000000000000",
16001 => "000000000000000000000000",
16002 => "000000000000000000000000",
16003 => "000000000000000000000000",
16004 => "000000000000000000000000",
16005 => "000000000000000000000000",
16006 => "000000000000000000000000",
16007 => "000000000000000000000000",
16008 => "000000000000000000000000",
16009 => "000000000000000000000000",
16010 => "000000000000000000000000",
16011 => "000000000000000000000000",
16012 => "000000000000000000000000",
16013 => "000000000000000000000000",
16014 => "000000000000000000000000",
16015 => "000000000000000000000000",
16016 => "000000000000000000000000",
16017 => "000000000000000000000000",
16018 => "000000000000000000000000",
16019 => "000111110001111100011111",
16020 => "010000110100001101000011",
16021 => "010000110100001101000011",
16022 => "010000110100001101000011",
16023 => "010000110100001101000011",
16024 => "000010110000101100001011",
16025 => "000000000000000000000000",
16026 => "000000000000000000000000",
16027 => "000000000000000000000000",
16028 => "000000000000000000000000",
16029 => "000000000000000000000000",
16030 => "000000000000000000000000",
16031 => "000000000000000000000000",
16032 => "000000000000000000000000",
16033 => "000000000000000000000000",
16034 => "000000000000000000000000",
16035 => "000000000000000000000000",
16036 => "000000000000000000000000",
16037 => "000000000000000000000000",
16038 => "000000000000000000000000",
16039 => "000000000000000000000000",
16040 => "000000000000000000000000",
16041 => "000000000000000000000000",
16042 => "000000000000000000000000",
16043 => "000000000000000000000000",
16044 => "000000000000000000000000",
16045 => "000000000000000000000000",
16046 => "000000000000000000000000",
16047 => "000000000000000000000000",
16048 => "000000000000000000000000",
16049 => "000000000000000000000000",
16050 => "000000000000000000000000",
16051 => "000000000000000000000000",
16052 => "000000000000000000000000",
16053 => "000000000000000000000000",
16054 => "000000000000000000000000",
16055 => "000000000000000000000000",
16056 => "000000000000000000000000",
16057 => "000000000000000000000000",
16058 => "000000000000000000000000",
16059 => "000000000000000000000000",
16060 => "000000000000000000000000",
16061 => "000000000000000000000000",
16062 => "000000000000000000000000",
16063 => "000000000000000000000000",
16064 => "001101100011011000110110",
16065 => "001101100011011000110110",
16066 => "001101100011011000110110",
16067 => "001101100011011000110110",
16068 => "001010010010100100101001",
16069 => "000000000000000000000000",
16070 => "000000000000000000000000",
16071 => "000000000000000000000000",
16072 => "000000000000000000000000",
16073 => "000000000000000000000000",
16074 => "000000000000000000000000",
16075 => "000000000000000000000000",
16076 => "000000000000000000000000",
16077 => "000000000000000000000000",
16078 => "000000000000000000000000",
16079 => "000000000000000000000000",
16080 => "000000000000000000000000",
16081 => "000000000000000000000000",
16082 => "000000000000000000000000",
16083 => "000000000000000000000000",
16084 => "000000000000000000000000",
16085 => "000000000000000000000000",
16086 => "000000000000000000000000",
16087 => "000000000000000000000000",
16088 => "000000000000000000000000",
16089 => "000000000000000000000000",
16090 => "000000000000000000000000",
16091 => "000000000000000000000000",
16092 => "000000000000000000000000",
16093 => "000000000000000000000000",
16094 => "000000000000000000000000",
16095 => "000000000000000000000000",
16096 => "000000000000000000000000",
16097 => "000000000000000000000000",
16098 => "000000000000000000000000",
16099 => "000000000000000000000000",
16100 => "000000000000000000000000",
16101 => "000000000000000000000000",
16102 => "000000000000000000000000",
16103 => "000000000000000000000000",
16104 => "000000000000000000000000",
16105 => "000000000000000000000000",
16106 => "010100000101000001010000",
16107 => "011001100110011001100110",
16108 => "010110000101100001011000",
16109 => "010000110100001101000011",
16110 => "010000110100001101000011",
16111 => "010000110100001101000011",
16112 => "010000110100001101000011",
16113 => "010000110100001101000011",
16114 => "010000110100001101000011",
16115 => "010100000101000001010000",
16116 => "011001100110011001100110",
16117 => "011001010110010101100101",
16118 => "010000110100001101000011",
16119 => "010000110100001101000011",
16120 => "010110110101101101011011",
16121 => "011001100110011001100110",
16122 => "010110100101101001011010",
16123 => "010000110100001101000011",
16124 => "010000110100001101000011",
16125 => "010000110100001101000011",
16126 => "010000110100001101000011",
16127 => "010000110100001101000011",
16128 => "010000110100001101000011",
16129 => "010011100100111001001110",
16130 => "011001100110011001100110",
16131 => "011001100110011001100110",
16132 => "000000000000000000000000",
16133 => "000000000000000000000000",
16134 => "000000000000000000000000",
16135 => "000000000000000000000000",
16136 => "000000000000000000000000",
16137 => "000000000000000000000000",
16138 => "000000000000000000000000",
16139 => "000000000000000000000000",
16140 => "000000000000000000000000",
16141 => "000000000000000000000000",
16142 => "000000000000000000000000",
16143 => "000000000000000000000000",
16144 => "000000000000000000000000",
16145 => "000000000000000000000000",
16146 => "000000000000000000000000",
16147 => "000000000000000000000000",
16148 => "000000000000000000000000",
16149 => "000000000000000000000000",
16150 => "000000000000000000000000",
16151 => "000000000000000000000000",
16152 => "000000000000000000000000",
16153 => "000000000000000000000000",
16154 => "000000000000000000000000",
16155 => "000000000000000000000000",
16156 => "000000000000000000000000",
16157 => "000000000000000000000000",
16158 => "000000000000000000000000",
16159 => "000000000000000000000000",
16160 => "000000000000000000000000",
16161 => "000000000000000000000000",
16162 => "000000000000000000000000",
16163 => "000000000000000000000000",
16164 => "000000000000000000000000",
16165 => "000000000000000000000000",
16166 => "000000000000000000000000",
16167 => "000000000000000000000000",
16168 => "000000000000000000000000",
16169 => "000110100001101000011010",
16170 => "001101100011011000110110",
16171 => "001101100011011000110110",
16172 => "001101100011011000110110",
16173 => "001101100011011000110110",
16174 => "000010010000100100001001",
16175 => "000000000000000000000000",
16176 => "000000000000000000000000",
16177 => "000000000000000000000000",
16178 => "000000000000000000000000",
16179 => "000000000000000000000000",
16180 => "000000000000000000000000",
16181 => "000000000000000000000000",
16182 => "000000000000000000000000",
16183 => "000000000000000000000000",
16184 => "000000000000000000000000",
16185 => "000000000000000000000000",
16186 => "000000000000000000000000",
16187 => "000000000000000000000000",
16188 => "000000000000000000000000",
16189 => "000000000000000000000000",
16190 => "000000000000000000000000",
16191 => "000000000000000000000000",
16192 => "000000000000000000000000",
16193 => "000000000000000000000000",
16194 => "000000000000000000000000",
16195 => "000000000000000000000000",
16196 => "000000000000000000000000",
16197 => "000000000000000000000000",
16198 => "000000000000000000000000",
16199 => "000000000000000000000000",
16200 => "000000000000000000000000",
16201 => "000000000000000000000000",
16202 => "000000000000000000000000",
16203 => "000000000000000000000000",
16204 => "000000000000000000000000",
16205 => "000000000000000000000000",
16206 => "000000000000000000000000",
16207 => "000000000000000000000000",
16208 => "000000000000000000000000",
16209 => "000000000000000000000000",
16210 => "000000000000000000000000",
16211 => "000000000000000000000000",
16212 => "000000000000000000000000",
16213 => "000000000000000000000000",
16214 => "000000000000000000000000",
16215 => "000000000000000000000000",
16216 => "000000000000000000000000",
16217 => "000000000000000000000000",
16218 => "000000000000000000000000",
16219 => "000000000000000000000000",
16220 => "000000000000000000000000",
16221 => "000000000000000000000000",
16222 => "000000000000000000000000",
16223 => "000000000000000000000000",
16224 => "000000000000000000000000",
16225 => "000000000000000000000000",
16226 => "000000000000000000000000",
16227 => "000000000000000000000000",
16228 => "000000000000000000000000",
16229 => "000000000000000000000000",
16230 => "000000000000000000000000",
16231 => "000000000000000000000000",
16232 => "000000000000000000000000",
16233 => "000000000000000000000000",
16234 => "000000000000000000000000",
16235 => "000000000000000000000000",
16236 => "000000000000000000000000",
16237 => "000000000000000000000000",
16238 => "000000000000000000000000",
16239 => "000000000000000000000000",
16240 => "000000000000000000000000",
16241 => "000000000000000000000000",
16242 => "000000000000000000000000",
16243 => "000000000000000000000000",
16244 => "000000000000000000000000",
16245 => "000000000000000000000000",
16246 => "000000000000000000000000",
16247 => "000000000000000000000000",
16248 => "000000000000000000000000",
16249 => "000000000000000000000000",
16250 => "000000000000000000000000",
16251 => "000000000000000000000000",
16252 => "000000000000000000000000",
16253 => "000000000000000000000000",
16254 => "000000000000000000000000",
16255 => "000000000000000000000000",
16256 => "010100000101000001010000",
16257 => "011001100110011001100110",
16258 => "010110000101100001011000",
16259 => "010000110100001101000011",
16260 => "010000110100001101000011",
16261 => "010000110100001101000011",
16262 => "010000110100001101000011",
16263 => "010000110100001101000011",
16264 => "010000110100001101000011",
16265 => "010100000101000001010000",
16266 => "011001100110011001100110",
16267 => "011001010110010101100101",
16268 => "010000110100001101000011",
16269 => "010000110100001101000011",
16270 => "010110110101101101011011",
16271 => "011001100110011001100110",
16272 => "010110100101101001011010",
16273 => "010000110100001101000011",
16274 => "010000110100001101000011",
16275 => "010000110100001101000011",
16276 => "010000110100001101000011",
16277 => "010000110100001101000011",
16278 => "010000110100001101000011",
16279 => "010011100100111001001110",
16280 => "011001100110011001100110",
16281 => "011001100110011001100110",
16282 => "000000000000000000000000",
16283 => "000000000000000000000000",
16284 => "000000000000000000000000",
16285 => "000000000000000000000000",
16286 => "000000000000000000000000",
16287 => "000000000000000000000000",
16288 => "000000000000000000000000",
16289 => "000000000000000000000000",
16290 => "000000000000000000000000",
16291 => "000000000000000000000000",
16292 => "000000000000000000000000",
16293 => "000000000000000000000000",
16294 => "000000000000000000000000",
16295 => "000000000000000000000000",
16296 => "000000000000000000000000",
16297 => "000000000000000000000000",
16298 => "000000000000000000000000",
16299 => "000000000000000000000000",
16300 => "000000000000000000000000",
16301 => "000000000000000000000000",
16302 => "000000000000000000000000",
16303 => "000000000000000000000000",
16304 => "000000000000000000000000",
16305 => "000000000000000000000000",
16306 => "000000000000000000000000",
16307 => "000000000000000000000000",
16308 => "000000000000000000000000",
16309 => "000000000000000000000000",
16310 => "000000000000000000000000",
16311 => "000000000000000000000000",
16312 => "000000000000000000000000",
16313 => "000000000000000000000000",
16314 => "000000000000000000000000",
16315 => "000000000000000000000000",
16316 => "000000000000000000000000",
16317 => "000000000000000000000000",
16318 => "000000000000000000000000",
16319 => "000000000000000000000000",
16320 => "000000000000000000000000",
16321 => "000000000000000000000000",
16322 => "000000000000000000000000",
16323 => "000000000000000000000000",
16324 => "000000000000000000000000",
16325 => "000000000000000000000000",
16326 => "000000000000000000000000",
16327 => "000000000000000000000000",
16328 => "000000000000000000000000",
16329 => "000000000000000000000000",
16330 => "000000000000000000000000",
16331 => "000000000000000000000000",
16332 => "000000000000000000000000",
16333 => "000000000000000000000000",
16334 => "000000000000000000000000",
16335 => "000000000000000000000000",
16336 => "000000000000000000000000",
16337 => "000000000000000000000000",
16338 => "000000000000000000000000",
16339 => "000000000000000000000000",
16340 => "000000000000000000000000",
16341 => "000000000000000000000000",
16342 => "000000000000000000000000",
16343 => "000000000000000000000000",
16344 => "000000000000000000000000",
16345 => "000000000000000000000000",
16346 => "000000000000000000000000",
16347 => "000000000000000000000000",
16348 => "000000000000000000000000",
16349 => "000000000000000000000000",
16350 => "000000000000000000000000",
16351 => "000000000000000000000000",
16352 => "000000000000000000000000",
16353 => "000000000000000000000000",
16354 => "000000000000000000000000",
16355 => "000000000000000000000000",
16356 => "000000000000000000000000",
16357 => "000000000000000000000000",
16358 => "000000000000000000000000",
16359 => "000000000000000000000000",
16360 => "000000000000000000000000",
16361 => "000000000000000000000000",
16362 => "000000000000000000000000",
16363 => "000000000000000000000000",
16364 => "000000000000000000000000",
16365 => "000000000000000000000000",
16366 => "000000000000000000000000",
16367 => "000000000000000000000000",
16368 => "000000000000000000000000",
16369 => "000000000000000000000000",
16370 => "000000000000000000000000",
16371 => "000000000000000000000000",
16372 => "000000000000000000000000",
16373 => "000000000000000000000000",
16374 => "000000000000000000000000",
16375 => "000000000000000000000000",
16376 => "000000000000000000000000",
16377 => "000000000000000000000000",
16378 => "000000000000000000000000",
16379 => "000000000000000000000000",
16380 => "000000000000000000000000",
16381 => "000000000000000000000000",
16382 => "000000000000000000000000",
16383 => "000000000000000000000000",
16384 => "000000000000000000000000",
16385 => "000000000000000000000000",
16386 => "000000000000000000000000",
16387 => "000000000000000000000000",
16388 => "000000000000000000000000",
16389 => "000000000000000000000000",
16390 => "000000000000000000000000",
16391 => "000000000000000000000000",
16392 => "000000000000000000000000",
16393 => "000000000000000000000000",
16394 => "000000000000000000000000",
16395 => "000000000000000000000000",
16396 => "000000000000000000000000",
16397 => "000000000000000000000000",
16398 => "000000000000000000000000",
16399 => "000000000000000000000000",
16400 => "000000000000000000000000",
16401 => "000000000000000000000000",
16402 => "000000000000000000000000",
16403 => "000000000000000000000000",
16404 => "000000000000000000000000",
16405 => "000000000000000000000000",
16406 => "010100000101000001010000",
16407 => "011001100110011001100110",
16408 => "010110000101100001011000",
16409 => "010000110100001101000011",
16410 => "010000110100001101000011",
16411 => "010000110100001101000011",
16412 => "010000110100001101000011",
16413 => "010000110100001101000011",
16414 => "010000110100001101000011",
16415 => "010100000101000001010000",
16416 => "011001100110011001100110",
16417 => "011001010110010101100101",
16418 => "010000110100001101000011",
16419 => "010000110100001101000011",
16420 => "010110110101101101011011",
16421 => "011001100110011001100110",
16422 => "010110100101101001011010",
16423 => "010000110100001101000011",
16424 => "010000110100001101000011",
16425 => "010000110100001101000011",
16426 => "010000110100001101000011",
16427 => "010000110100001101000011",
16428 => "010000110100001101000011",
16429 => "010011100100111001001110",
16430 => "011001100110011001100110",
16431 => "011001100110011001100110",
16432 => "000000000000000000000000",
16433 => "000000000000000000000000",
16434 => "000000000000000000000000",
16435 => "000000000000000000000000",
16436 => "000000000000000000000000",
16437 => "000000000000000000000000",
16438 => "000000000000000000000000",
16439 => "000000000000000000000000",
16440 => "000000000000000000000000",
16441 => "000000000000000000000000",
16442 => "000000000000000000000000",
16443 => "000000000000000000000000",
16444 => "000000000000000000000000",
16445 => "000000000000000000000000",
16446 => "000000000000000000000000",
16447 => "000000000000000000000000",
16448 => "000000000000000000000000",
16449 => "000000000000000000000000",
16450 => "000000000000000000000000",
16451 => "000000000000000000000000",
16452 => "000000000000000000000000",
16453 => "000000000000000000000000",
16454 => "000000000000000000000000",
16455 => "000000000000000000000000",
16456 => "000000000000000000000000",
16457 => "000000000000000000000000",
16458 => "000000000000000000000000",
16459 => "000000000000000000000000",
16460 => "000000000000000000000000",
16461 => "000000000000000000000000",
16462 => "000000000000000000000000",
16463 => "000000000000000000000000",
16464 => "000000000000000000000000",
16465 => "000000000000000000000000",
16466 => "000000000000000000000000",
16467 => "000000000000000000000000",
16468 => "000000000000000000000000",
16469 => "000000000000000000000000",
16470 => "000000000000000000000000",
16471 => "000000000000000000000000",
16472 => "000000000000000000000000",
16473 => "000000000000000000000000",
16474 => "000000000000000000000000",
16475 => "000000000000000000000000",
16476 => "000000000000000000000000",
16477 => "000000000000000000000000",
16478 => "000000000000000000000000",
16479 => "000000000000000000000000",
16480 => "000000000000000000000000",
16481 => "000000000000000000000000",
16482 => "000000000000000000000000",
16483 => "000000000000000000000000",
16484 => "000000000000000000000000",
16485 => "000000000000000000000000",
16486 => "000000000000000000000000",
16487 => "000000000000000000000000",
16488 => "000000000000000000000000",
16489 => "000000000000000000000000",
16490 => "000000000000000000000000",
16491 => "000000000000000000000000",
16492 => "000000000000000000000000",
16493 => "000000000000000000000000",
16494 => "000000000000000000000000",
16495 => "000000000000000000000000",
16496 => "000000000000000000000000",
16497 => "000000000000000000000000",
16498 => "000000000000000000000000",
16499 => "000000000000000000000000",
16500 => "000000000000000000000000",
16501 => "000000000000000000000000",
16502 => "000000000000000000000000",
16503 => "000000000000000000000000",
16504 => "000000000000000000000000",
16505 => "000000000000000000000000",
16506 => "000000000000000000000000",
16507 => "000000000000000000000000",
16508 => "000000000000000000000000",
16509 => "000000000000000000000000",
16510 => "000000000000000000000000",
16511 => "000000000000000000000000",
16512 => "000000000000000000000000",
16513 => "000000000000000000000000",
16514 => "000000000000000000000000",
16515 => "000000000000000000000000",
16516 => "000000000000000000000000",
16517 => "000000000000000000000000",
16518 => "000000000000000000000000",
16519 => "000000000000000000000000",
16520 => "000000000000000000000000",
16521 => "000000000000000000000000",
16522 => "000000000000000000000000",
16523 => "000000000000000000000000",
16524 => "000000000000000000000000",
16525 => "000000000000000000000000",
16526 => "000000000000000000000000",
16527 => "000000000000000000000000",
16528 => "000000000000000000000000",
16529 => "000000000000000000000000",
16530 => "000000000000000000000000",
16531 => "000000000000000000000000",
16532 => "000000000000000000000000",
16533 => "000000000000000000000000",
16534 => "000000000000000000000000",
16535 => "000000000000000000000000",
16536 => "000000000000000000000000",
16537 => "000000000000000000000000",
16538 => "000000000000000000000000",
16539 => "000000000000000000000000",
16540 => "000000000000000000000000",
16541 => "000000000000000000000000",
16542 => "000000000000000000000000",
16543 => "000000000000000000000000",
16544 => "000000000000000000000000",
16545 => "000000000000000000000000",
16546 => "000000000000000000000000",
16547 => "000000000000000000000000",
16548 => "000000000000000000000000",
16549 => "000000000000000000000000",
16550 => "000000000000000000000000",
16551 => "000000000000000000000000",
16552 => "000000000000000000000000",
16553 => "000000000000000000000000",
16554 => "000000000000000000000000",
16555 => "000000000000000000000000",
16556 => "010100000101000001010000",
16557 => "011001100110011001100110",
16558 => "010110000101100001011000",
16559 => "010000110100001101000011",
16560 => "010000110100001101000011",
16561 => "010000110100001101000011",
16562 => "010000110100001101000011",
16563 => "010000110100001101000011",
16564 => "010000110100001101000011",
16565 => "010100000101000001010000",
16566 => "011001100110011001100110",
16567 => "011001010110010101100101",
16568 => "010000110100001101000011",
16569 => "010000110100001101000011",
16570 => "010110110101101101011011",
16571 => "011001100110011001100110",
16572 => "010110100101101001011010",
16573 => "010000110100001101000011",
16574 => "010000110100001101000011",
16575 => "010000110100001101000011",
16576 => "010000110100001101000011",
16577 => "010000110100001101000011",
16578 => "010000110100001101000011",
16579 => "010011100100111001001110",
16580 => "011001100110011001100110",
16581 => "011001100110011001100110",
16582 => "000000000000000000000000",
16583 => "000000000000000000000000",
16584 => "000000000000000000000000",
16585 => "000000000000000000000000",
16586 => "000000000000000000000000",
16587 => "000000000000000000000000",
16588 => "000000000000000000000000",
16589 => "000000000000000000000000",
16590 => "000000000000000000000000",
16591 => "000000000000000000000000",
16592 => "000000000000000000000000",
16593 => "000000000000000000000000",
16594 => "000000000000000000000000",
16595 => "000000000000000000000000",
16596 => "000000000000000000000000",
16597 => "000000000000000000000000",
16598 => "000000000000000000000000",
16599 => "000000000000000000000000",
16600 => "000000000000000000000000",
16601 => "000000000000000000000000",
16602 => "000000000000000000000000",
16603 => "000000000000000000000000",
16604 => "000000000000000000000000",
16605 => "000000000000000000000000",
16606 => "000000000000000000000000",
16607 => "000000000000000000000000",
16608 => "000000000000000000000000",
16609 => "000000000000000000000000",
16610 => "000000000000000000000000",
16611 => "000000000000000000000000",
16612 => "000000000000000000000000",
16613 => "000000000000000000000000",
16614 => "000000000000000000000000",
16615 => "000000000000000000000000",
16616 => "000000000000000000000000",
16617 => "000000000000000000000000",
16618 => "000000000000000000000000",
16619 => "000000000000000000000000",
16620 => "000000000000000000000000",
16621 => "000000000000000000000000",
16622 => "000000000000000000000000",
16623 => "000000000000000000000000",
16624 => "000000000000000000000000",
16625 => "000000000000000000000000",
16626 => "000000000000000000000000",
16627 => "000000000000000000000000",
16628 => "000000000000000000000000",
16629 => "000000000000000000000000",
16630 => "000000000000000000000000",
16631 => "000000000000000000000000",
16632 => "000000000000000000000000",
16633 => "000000000000000000000000",
16634 => "000000000000000000000000",
16635 => "000000000000000000000000",
16636 => "000000000000000000000000",
16637 => "000000000000000000000000",
16638 => "000000000000000000000000",
16639 => "000000000000000000000000",
16640 => "000000000000000000000000",
16641 => "000000000000000000000000",
16642 => "000000000000000000000000",
16643 => "000000000000000000000000",
16644 => "000000000000000000000000",
16645 => "000000000000000000000000",
16646 => "000000000000000000000000",
16647 => "000000000000000000000000",
16648 => "000000000000000000000000",
16649 => "000000000000000000000000",
16650 => "000000000000000000000000",
16651 => "000000000000000000000000",
16652 => "000000000000000000000000",
16653 => "000000000000000000000000",
16654 => "000000000000000000000000",
16655 => "000000000000000000000000",
16656 => "000000000000000000000000",
16657 => "000000000000000000000000",
16658 => "000000000000000000000000",
16659 => "000000000000000000000000",
16660 => "000000000000000000000000",
16661 => "000000000000000000000000",
16662 => "000000000000000000000000",
16663 => "000000000000000000000000",
16664 => "000000000000000000000000",
16665 => "000000000000000000000000",
16666 => "000000000000000000000000",
16667 => "000000000000000000000000",
16668 => "000000000000000000000000",
16669 => "000000000000000000000000",
16670 => "000000000000000000000000",
16671 => "000000000000000000000000",
16672 => "000000000000000000000000",
16673 => "000000000000000000000000",
16674 => "000000000000000000000000",
16675 => "000000000000000000000000",
16676 => "000000000000000000000000",
16677 => "000000000000000000000000",
16678 => "000000000000000000000000",
16679 => "000000000000000000000000",
16680 => "000000000000000000000000",
16681 => "000000000000000000000000",
16682 => "000000000000000000000000",
16683 => "000000000000000000000000",
16684 => "000000000000000000000000",
16685 => "000000000000000000000000",
16686 => "000000000000000000000000",
16687 => "000000000000000000000000",
16688 => "000000000000000000000000",
16689 => "000000000000000000000000",
16690 => "000000000000000000000000",
16691 => "000000000000000000000000",
16692 => "000000000000000000000000",
16693 => "000000000000000000000000",
16694 => "000000000000000000000000",
16695 => "000000000000000000000000",
16696 => "000000000000000000000000",
16697 => "000000000000000000000000",
16698 => "000000000000000000000000",
16699 => "000000000000000000000000",
16700 => "000000000000000000000000",
16701 => "000000000000000000000000",
16702 => "000000000000000000000000",
16703 => "000000000000000000000000",
16704 => "000000000000000000000000",
16705 => "000000000000000000000000",
16706 => "010100000101000001010000",
16707 => "011001100110011001100110",
16708 => "010110000101100001011000",
16709 => "010000110100001101000011",
16710 => "010000110100001101000011",
16711 => "010000110100001101000011",
16712 => "010000110100001101000011",
16713 => "010000110100001101000011",
16714 => "010000110100001101000011",
16715 => "010100000101000001010000",
16716 => "011001100110011001100110",
16717 => "011001010110010101100101",
16718 => "010000110100001101000011",
16719 => "010000110100001101000011",
16720 => "010110110101101101011011",
16721 => "011001100110011001100110",
16722 => "010110100101101001011010",
16723 => "010000110100001101000011",
16724 => "010000110100001101000011",
16725 => "010000110100001101000011",
16726 => "010000110100001101000011",
16727 => "010000110100001101000011",
16728 => "010000110100001101000011",
16729 => "010011100100111001001110",
16730 => "011001100110011001100110",
16731 => "011001100110011001100110",
16732 => "000000000000000000000000",
16733 => "000000000000000000000000",
16734 => "000000000000000000000000",
16735 => "000000000000000000000000",
16736 => "000000000000000000000000",
16737 => "000000000000000000000000",
16738 => "000000000000000000000000",
16739 => "000000000000000000000000",
16740 => "000000000000000000000000",
16741 => "000000000000000000000000",
16742 => "000000000000000000000000",
16743 => "000000000000000000000000",
16744 => "000000000000000000000000",
16745 => "000000000000000000000000",
16746 => "000000000000000000000000",
16747 => "000000000000000000000000",
16748 => "000000000000000000000000",
16749 => "000000000000000000000000",
16750 => "000000000000000000000000",
16751 => "000000000000000000000000",
16752 => "000000000000000000000000",
16753 => "000000000000000000000000",
16754 => "000000000000000000000000",
16755 => "000000000000000000000000",
16756 => "000000000000000000000000",
16757 => "000000000000000000000000",
16758 => "000000000000000000000000",
16759 => "000000000000000000000000",
16760 => "000000000000000000000000",
16761 => "000000000000000000000000",
16762 => "000000000000000000000000",
16763 => "000000000000000000000000",
16764 => "000000000000000000000000",
16765 => "000000000000000000000000",
16766 => "000000000000000000000000",
16767 => "000000000000000000000000",
16768 => "000000000000000000000000",
16769 => "000000000000000000000000",
16770 => "000000000000000000000000",
16771 => "000000000000000000000000",
16772 => "000000000000000000000000",
16773 => "000000000000000000000000",
16774 => "000000000000000000000000",
16775 => "000000000000000000000000",
16776 => "000000000000000000000000",
16777 => "000000000000000000000000",
16778 => "000000000000000000000000",
16779 => "000000000000000000000000",
16780 => "000000000000000000000000",
16781 => "000000000000000000000000",
16782 => "000000000000000000000000",
16783 => "000000000000000000000000",
16784 => "000000000000000000000000",
16785 => "000000000000000000000000",
16786 => "000000000000000000000000",
16787 => "000000000000000000000000",
16788 => "000000000000000000000000",
16789 => "000000000000000000000000",
16790 => "000000000000000000000000",
16791 => "000000000000000000000000",
16792 => "000000000000000000000000",
16793 => "000000000000000000000000",
16794 => "000000000000000000000000",
16795 => "000000000000000000000000",
16796 => "000000000000000000000000",
16797 => "000000000000000000000000",
16798 => "000000000000000000000000",
16799 => "000000000000000000000000",
16800 => "000000000000000000000000",
16801 => "000000000000000000000000",
16802 => "000000000000000000000000",
16803 => "000000000000000000000000",
16804 => "000000000000000000000000",
16805 => "000000000000000000000000",
16806 => "000000000000000000000000",
16807 => "000000000000000000000000",
16808 => "000000000000000000000000",
16809 => "000000000000000000000000",
16810 => "000000000000000000000000",
16811 => "000000000000000000000000",
16812 => "000000000000000000000000",
16813 => "000000000000000000000000",
16814 => "000000000000000000000000",
16815 => "000000000000000000000000",
16816 => "000000000000000000000000",
16817 => "000000000000000000000000",
16818 => "000000000000000000000000",
16819 => "000000000000000000000000",
16820 => "000000000000000000000000",
16821 => "000000000000000000000000",
16822 => "000000000000000000000000",
16823 => "000000000000000000000000",
16824 => "000000000000000000000000",
16825 => "000000000000000000000000",
16826 => "000000000000000000000000",
16827 => "000000000000000000000000",
16828 => "000000000000000000000000",
16829 => "000000000000000000000000",
16830 => "000000000000000000000000",
16831 => "000000000000000000000000",
16832 => "000000000000000000000000",
16833 => "000000000000000000000000",
16834 => "000000000000000000000000",
16835 => "000000000000000000000000",
16836 => "000000000000000000000000",
16837 => "000000000000000000000000",
16838 => "000000000000000000000000",
16839 => "000000000000000000000000",
16840 => "000000000000000000000000",
16841 => "000000000000000000000000",
16842 => "000000000000000000000000",
16843 => "000000000000000000000000",
16844 => "000000000000000000000000",
16845 => "000000000000000000000000",
16846 => "000000000000000000000000",
16847 => "000000000000000000000000",
16848 => "000000000000000000000000",
16849 => "000000000000000000000000",
16850 => "000000000000000000000000",
16851 => "000000000000000000000000",
16852 => "000000000000000000000000",
16853 => "000000110000001100000011",
16854 => "001000100010001000100010",
16855 => "001000100010001000100010",
16856 => "010101110101011101010111",
16857 => "011001100110011001100110",
16858 => "010110000101100001011000",
16859 => "010000110100001101000011",
16860 => "010000110100001101000011",
16861 => "010000110100001101000011",
16862 => "010000110100001101000011",
16863 => "010000110100001101000011",
16864 => "010000110100001101000011",
16865 => "010100000101000001010000",
16866 => "011001100110011001100110",
16867 => "011001010110010101100101",
16868 => "010000110100001101000011",
16869 => "010000110100001101000011",
16870 => "010110110101101101011011",
16871 => "011001100110011001100110",
16872 => "010110100101101001011010",
16873 => "010000110100001101000011",
16874 => "010000110100001101000011",
16875 => "010000110100001101000011",
16876 => "010000110100001101000011",
16877 => "010000110100001101000011",
16878 => "010000110100001101000011",
16879 => "010011100100111001001110",
16880 => "011001100110011001100110",
16881 => "011001100110011001100110",
16882 => "001000100010001000100010",
16883 => "001000100010001000100010",
16884 => "000011010000110100001101",
16885 => "000000000000000000000000",
16886 => "000000000000000000000000",
16887 => "000000000000000000000000",
16888 => "000000000000000000000000",
16889 => "000000000000000000000000",
16890 => "000000000000000000000000",
16891 => "000000000000000000000000",
16892 => "000000000000000000000000",
16893 => "000000000000000000000000",
16894 => "000000000000000000000000",
16895 => "000000000000000000000000",
16896 => "000000000000000000000000",
16897 => "000000000000000000000000",
16898 => "000000000000000000000000",
16899 => "000000000000000000000000",
16900 => "000000000000000000000000",
16901 => "000000000000000000000000",
16902 => "000000000000000000000000",
16903 => "000000000000000000000000",
16904 => "000000000000000000000000",
16905 => "000000000000000000000000",
16906 => "000000000000000000000000",
16907 => "000000000000000000000000",
16908 => "000000000000000000000000",
16909 => "000000000000000000000000",
16910 => "000000000000000000000000",
16911 => "000000000000000000000000",
16912 => "000000000000000000000000",
16913 => "000000000000000000000000",
16914 => "000000000000000000000000",
16915 => "000000000000000000000000",
16916 => "000000000000000000000000",
16917 => "000000000000000000000000",
16918 => "000000000000000000000000",
16919 => "000000000000000000000000",
16920 => "000000000000000000000000",
16921 => "000000000000000000000000",
16922 => "000000000000000000000000",
16923 => "000000000000000000000000",
16924 => "000000000000000000000000",
16925 => "000000000000000000000000",
16926 => "000000000000000000000000",
16927 => "000000000000000000000000",
16928 => "000000000000000000000000",
16929 => "000000000000000000000000",
16930 => "000000000000000000000000",
16931 => "000000000000000000000000",
16932 => "000000000000000000000000",
16933 => "000000000000000000000000",
16934 => "000000000000000000000000",
16935 => "000000000000000000000000",
16936 => "000000000000000000000000",
16937 => "000000000000000000000000",
16938 => "000000000000000000000000",
16939 => "000000000000000000000000",
16940 => "000000000000000000000000",
16941 => "000000000000000000000000",
16942 => "000000000000000000000000",
16943 => "000000000000000000000000",
16944 => "000000000000000000000000",
16945 => "000000000000000000000000",
16946 => "000000000000000000000000",
16947 => "000000000000000000000000",
16948 => "000000000000000000000000",
16949 => "000000000000000000000000",
16950 => "000000000000000000000000",
16951 => "000000000000000000000000",
16952 => "000000000000000000000000",
16953 => "000000000000000000000000",
16954 => "000000000000000000000000",
16955 => "000000000000000000000000",
16956 => "000000000000000000000000",
16957 => "000000000000000000000000",
16958 => "000000000000000000000000",
16959 => "000000000000000000000000",
16960 => "000000000000000000000000",
16961 => "000000000000000000000000",
16962 => "000000000000000000000000",
16963 => "000000000000000000000000",
16964 => "000000000000000000000000",
16965 => "000000000000000000000000",
16966 => "000000000000000000000000",
16967 => "000000000000000000000000",
16968 => "000000000000000000000000",
16969 => "000000000000000000000000",
16970 => "000000000000000000000000",
16971 => "000000000000000000000000",
16972 => "000000000000000000000000",
16973 => "000000000000000000000000",
16974 => "000000000000000000000000",
16975 => "000000000000000000000000",
16976 => "000000000000000000000000",
16977 => "000000000000000000000000",
16978 => "000000000000000000000000",
16979 => "000000000000000000000000",
16980 => "000000000000000000000000",
16981 => "000000000000000000000000",
16982 => "000000000000000000000000",
16983 => "000000000000000000000000",
16984 => "000000000000000000000000",
16985 => "000000000000000000000000",
16986 => "000000000000000000000000",
16987 => "000000000000000000000000",
16988 => "000000000000000000000000",
16989 => "000000000000000000000000",
16990 => "000000000000000000000000",
16991 => "000000000000000000000000",
16992 => "000000000000000000000000",
16993 => "000000000000000000000000",
16994 => "000000000000000000000000",
16995 => "000000000000000000000000",
16996 => "000000000000000000000000",
16997 => "000000000000000000000000",
16998 => "000000000000000000000000",
16999 => "000000000000000000000000",
17000 => "000000000000000000000000",
17001 => "000000000000000000000000",
17002 => "000000000000000000000000",
17003 => "000001100000011000000110",
17004 => "010000110100001101000011",
17005 => "010000110100001101000011",
17006 => "010111110101111101011111",
17007 => "011001100110011001100110",
17008 => "010110000101100001011000",
17009 => "010000110100001101000011",
17010 => "010000110100001101000011",
17011 => "010000110100001101000011",
17012 => "010000110100001101000011",
17013 => "010000110100001101000011",
17014 => "010000110100001101000011",
17015 => "010100000101000001010000",
17016 => "011001100110011001100110",
17017 => "011001010110010101100101",
17018 => "010000110100001101000011",
17019 => "010000110100001101000011",
17020 => "010110110101101101011011",
17021 => "011001100110011001100110",
17022 => "010110100101101001011010",
17023 => "010000110100001101000011",
17024 => "010000110100001101000011",
17025 => "010000110100001101000011",
17026 => "010000110100001101000011",
17027 => "010000110100001101000011",
17028 => "010000110100001101000011",
17029 => "010011100100111001001110",
17030 => "011001100110011001100110",
17031 => "011001100110011001100110",
17032 => "010000110100001101000011",
17033 => "010000110100001101000011",
17034 => "000110010001100100011001",
17035 => "000000000000000000000000",
17036 => "000000000000000000000000",
17037 => "000000000000000000000000",
17038 => "000000000000000000000000",
17039 => "000000000000000000000000",
17040 => "000000000000000000000000",
17041 => "000000000000000000000000",
17042 => "000000000000000000000000",
17043 => "000000000000000000000000",
17044 => "000000000000000000000000",
17045 => "000000000000000000000000",
17046 => "000000000000000000000000",
17047 => "000000000000000000000000",
17048 => "000000000000000000000000",
17049 => "000000000000000000000000",
17050 => "000000000000000000000000",
17051 => "000000000000000000000000",
17052 => "000000000000000000000000",
17053 => "000000000000000000000000",
17054 => "000000000000000000000000",
17055 => "000000000000000000000000",
17056 => "000000000000000000000000",
17057 => "000000000000000000000000",
17058 => "000000000000000000000000",
17059 => "000000000000000000000000",
17060 => "000000000000000000000000",
17061 => "000000000000000000000000",
17062 => "000000000000000000000000",
17063 => "000000000000000000000000",
17064 => "000000000000000000000000",
17065 => "000000000000000000000000",
17066 => "000000000000000000000000",
17067 => "000000000000000000000000",
17068 => "000000000000000000000000",
17069 => "000000000000000000000000",
17070 => "000000000000000000000000",
17071 => "000000000000000000000000",
17072 => "000000000000000000000000",
17073 => "000000000000000000000000",
17074 => "000000000000000000000000",
17075 => "000000000000000000000000",
17076 => "000000000000000000000000",
17077 => "000000000000000000000000",
17078 => "000000000000000000000000",
17079 => "000000000000000000000000",
17080 => "000000000000000000000000",
17081 => "000000000000000000000000",
17082 => "000000000000000000000000",
17083 => "000000000000000000000000",
17084 => "000000000000000000000000",
17085 => "000000000000000000000000",
17086 => "000000000000000000000000",
17087 => "000000000000000000000000",
17088 => "000000000000000000000000",
17089 => "000000000000000000000000",
17090 => "000000000000000000000000",
17091 => "000000000000000000000000",
17092 => "000000000000000000000000",
17093 => "000000000000000000000000",
17094 => "000000000000000000000000",
17095 => "000000000000000000000000",
17096 => "000000000000000000000000",
17097 => "000000000000000000000000",
17098 => "000000000000000000000000",
17099 => "000000000000000000000000",
17100 => "000000000000000000000000",
17101 => "000000000000000000000000",
17102 => "000000000000000000000000",
17103 => "000000000000000000000000",
17104 => "000000000000000000000000",
17105 => "000000000000000000000000",
17106 => "000000000000000000000000",
17107 => "000000000000000000000000",
17108 => "000000000000000000000000",
17109 => "000000000000000000000000",
17110 => "000000000000000000000000",
17111 => "000000000000000000000000",
17112 => "000000000000000000000000",
17113 => "000000000000000000000000",
17114 => "000000000000000000000000",
17115 => "000000000000000000000000",
17116 => "000000000000000000000000",
17117 => "000000000000000000000000",
17118 => "000000000000000000000000",
17119 => "000000000000000000000000",
17120 => "000000000000000000000000",
17121 => "000000000000000000000000",
17122 => "000000000000000000000000",
17123 => "000000000000000000000000",
17124 => "000000000000000000000000",
17125 => "000000000000000000000000",
17126 => "000000000000000000000000",
17127 => "000000000000000000000000",
17128 => "000000000000000000000000",
17129 => "000000000000000000000000",
17130 => "000000000000000000000000",
17131 => "000000000000000000000000",
17132 => "000000000000000000000000",
17133 => "000000000000000000000000",
17134 => "000000000000000000000000",
17135 => "000000000000000000000000",
17136 => "000000000000000000000000",
17137 => "000000000000000000000000",
17138 => "000000000000000000000000",
17139 => "000000000000000000000000",
17140 => "000000000000000000000000",
17141 => "000000000000000000000000",
17142 => "000000000000000000000000",
17143 => "000000000000000000000000",
17144 => "000000000000000000000000",
17145 => "000000000000000000000000",
17146 => "000000000000000000000000",
17147 => "000000000000000000000000",
17148 => "000000000000000000000000",
17149 => "000000000000000000000000",
17150 => "000000000000000000000000",
17151 => "000000000000000000000000",
17152 => "000000000000000000000000",
17153 => "000001110000011100000111",
17154 => "010010000100100001001000",
17155 => "010010000100100001001000",
17156 => "010110110101101101011011",
17157 => "011000010110000101100001",
17158 => "010101110101011101010111",
17159 => "010010000100100001001000",
17160 => "010010000100100001001000",
17161 => "010000110100001101000011",
17162 => "010000110100001101000011",
17163 => "010000110100001101000011",
17164 => "010000110100001101000011",
17165 => "010100000101000001010000",
17166 => "011001100110011001100110",
17167 => "011001010110010101100101",
17168 => "010000110100001101000011",
17169 => "010000110100001101000011",
17170 => "010110110101101101011011",
17171 => "011001100110011001100110",
17172 => "010110100101101001011010",
17173 => "010000110100001101000011",
17174 => "010000110100001101000011",
17175 => "010000110100001101000011",
17176 => "010000110100001101000011",
17177 => "010001110100011101000111",
17178 => "010010000100100001001000",
17179 => "010100000101000001010000",
17180 => "011000010110000101100001",
17181 => "011000010110000101100001",
17182 => "010010010100100101001001",
17183 => "010010000100100001001000",
17184 => "000110110001101100011011",
17185 => "000000000000000000000000",
17186 => "000000000000000000000000",
17187 => "000000000000000000000000",
17188 => "000000000000000000000000",
17189 => "000000000000000000000000",
17190 => "000000000000000000000000",
17191 => "000000000000000000000000",
17192 => "000000000000000000000000",
17193 => "000000000000000000000000",
17194 => "000000000000000000000000",
17195 => "000000000000000000000000",
17196 => "000000000000000000000000",
17197 => "000000000000000000000000",
17198 => "000000000000000000000000",
17199 => "000000000000000000000000",
17200 => "000000000000000000000000",
17201 => "000000000000000000000000",
17202 => "000000000000000000000000",
17203 => "000000000000000000000000",
17204 => "000000000000000000000000",
17205 => "000000000000000000000000",
17206 => "000000000000000000000000",
17207 => "000000000000000000000000",
17208 => "000000000000000000000000",
17209 => "000000000000000000000000",
17210 => "000000000000000000000000",
17211 => "000000000000000000000000",
17212 => "000000000000000000000000",
17213 => "000000000000000000000000",
17214 => "000000000000000000000000",
17215 => "000000000000000000000000",
17216 => "000000000000000000000000",
17217 => "000000000000000000000000",
17218 => "000000000000000000000000",
17219 => "000000000000000000000000",
17220 => "000000000000000000000000",
17221 => "000000000000000000000000",
17222 => "000000000000000000000000",
17223 => "000000000000000000000000",
17224 => "000000000000000000000000",
17225 => "000000000000000000000000",
17226 => "000000000000000000000000",
17227 => "000000000000000000000000",
17228 => "000000000000000000000000",
17229 => "000000000000000000000000",
17230 => "000000000000000000000000",
17231 => "000000000000000000000000",
17232 => "000000000000000000000000",
17233 => "000000000000000000000000",
17234 => "000000000000000000000000",
17235 => "000000000000000000000000",
17236 => "000000000000000000000000",
17237 => "000000000000000000000000",
17238 => "000000000000000000000000",
17239 => "000000000000000000000000",
17240 => "000000000000000000000000",
17241 => "000000000000000000000000",
17242 => "000000000000000000000000",
17243 => "000000000000000000000000",
17244 => "000000000000000000000000",
17245 => "000000000000000000000000",
17246 => "000000000000000000000000",
17247 => "000000000000000000000000",
17248 => "000000000000000000000000",
17249 => "000000000000000000000000",
17250 => "000000000000000000000000",
17251 => "000000000000000000000000",
17252 => "000000000000000000000000",
17253 => "000000000000000000000000",
17254 => "000000000000000000000000",
17255 => "000000000000000000000000",
17256 => "000000000000000000000000",
17257 => "000000000000000000000000",
17258 => "000000000000000000000000",
17259 => "000000000000000000000000",
17260 => "000000000000000000000000",
17261 => "000000000000000000000000",
17262 => "000000000000000000000000",
17263 => "000000000000000000000000",
17264 => "000000000000000000000000",
17265 => "000000000000000000000000",
17266 => "000000000000000000000000",
17267 => "000000000000000000000000",
17268 => "000000000000000000000000",
17269 => "000000000000000000000000",
17270 => "000000000000000000000000",
17271 => "000000000000000000000000",
17272 => "000000000000000000000000",
17273 => "000000000000000000000000",
17274 => "000000000000000000000000",
17275 => "000000000000000000000000",
17276 => "000000000000000000000000",
17277 => "000000000000000000000000",
17278 => "000000000000000000000000",
17279 => "000000000000000000000000",
17280 => "000000000000000000000000",
17281 => "000000000000000000000000",
17282 => "000000000000000000000000",
17283 => "000000000000000000000000",
17284 => "000000000000000000000000",
17285 => "000000000000000000000000",
17286 => "000000000000000000000000",
17287 => "000000000000000000000000",
17288 => "000000000000000000000000",
17289 => "000000000000000000000000",
17290 => "000000000000000000000000",
17291 => "000000000000000000000000",
17292 => "000000000000000000000000",
17293 => "000000000000000000000000",
17294 => "000000000000000000000000",
17295 => "000000000000000000000000",
17296 => "000000000000000000000000",
17297 => "000000000000000000000000",
17298 => "000000000000000000000000",
17299 => "000000000000000000000000",
17300 => "000000000000000000000000",
17301 => "000000000000000000000000",
17302 => "000000000000000000000000",
17303 => "000010100000101000001010",
17304 => "011001100110011001100110",
17305 => "011001100110011001100110",
17306 => "010010100100101001001010",
17307 => "010000110100001101000011",
17308 => "010100010101000101010001",
17309 => "011001100110011001100110",
17310 => "011001000110010001100100",
17311 => "010000110100001101000011",
17312 => "010000110100001101000011",
17313 => "010000110100001101000011",
17314 => "010000110100001101000011",
17315 => "010100000101000001010000",
17316 => "011001100110011001100110",
17317 => "011001010110010101100101",
17318 => "010000110100001101000011",
17319 => "010000110100001101000011",
17320 => "010110110101101101011011",
17321 => "011001100110011001100110",
17322 => "010110100101101001011010",
17323 => "010000110100001101000011",
17324 => "010000110100001101000011",
17325 => "010000110100001101000011",
17326 => "010000110100001101000011",
17327 => "010110100101101001011010",
17328 => "011001100110011001100110",
17329 => "010110110101101101011011",
17330 => "010000110100001101000011",
17331 => "010000110100001101000011",
17332 => "011001100110011001100110",
17333 => "011001100110011001100110",
17334 => "001001100010011000100110",
17335 => "000000000000000000000000",
17336 => "000000000000000000000000",
17337 => "000000000000000000000000",
17338 => "000000000000000000000000",
17339 => "000000000000000000000000",
17340 => "000000000000000000000000",
17341 => "000000000000000000000000",
17342 => "000000000000000000000000",
17343 => "000000000000000000000000",
17344 => "000000000000000000000000",
17345 => "000000000000000000000000",
17346 => "000000000000000000000000",
17347 => "000000000000000000000000",
17348 => "000000000000000000000000",
17349 => "000000000000000000000000",
17350 => "000000000000000000000000",
17351 => "000000000000000000000000",
17352 => "000000000000000000000000",
17353 => "000000000000000000000000",
17354 => "000000000000000000000000",
17355 => "000000000000000000000000",
17356 => "000000000000000000000000",
17357 => "000000000000000000000000",
17358 => "000000000000000000000000",
17359 => "000000000000000000000000",
17360 => "000000000000000000000000",
17361 => "000000000000000000000000",
17362 => "000000000000000000000000",
17363 => "000000000000000000000000",
17364 => "000000000000000000000000",
17365 => "000000000000000000000000",
17366 => "000000000000000000000000",
17367 => "000000000000000000000000",
17368 => "000000000000000000000000",
17369 => "000000000000000000000000",
17370 => "000000000000000000000000",
17371 => "000000000000000000000000",
17372 => "000000000000000000000000",
17373 => "000000000000000000000000",
17374 => "000000000000000000000000",
17375 => "000000000000000000000000",
17376 => "000000000000000000000000",
17377 => "000000000000000000000000",
17378 => "000000000000000000000000",
17379 => "000000000000000000000000",
17380 => "000000000000000000000000",
17381 => "000000000000000000000000",
17382 => "000000000000000000000000",
17383 => "000000000000000000000000",
17384 => "000000000000000000000000",
17385 => "000000000000000000000000",
17386 => "000000000000000000000000",
17387 => "000000000000000000000000",
17388 => "000000000000000000000000",
17389 => "000000000000000000000000",
17390 => "000000000000000000000000",
17391 => "000000000000000000000000",
17392 => "000000000000000000000000",
17393 => "000000000000000000000000",
17394 => "000000000000000000000000",
17395 => "000000000000000000000000",
17396 => "000000000000000000000000",
17397 => "000000000000000000000000",
17398 => "000000000000000000000000",
17399 => "000000000000000000000000",
17400 => "000000000000000000000000",
17401 => "000000000000000000000000",
17402 => "000000000000000000000000",
17403 => "000000000000000000000000",
17404 => "000000000000000000000000",
17405 => "000000000000000000000000",
17406 => "000000000000000000000000",
17407 => "000000000000000000000000",
17408 => "000000000000000000000000",
17409 => "000000000000000000000000",
17410 => "000000000000000000000000",
17411 => "000000000000000000000000",
17412 => "000000000000000000000000",
17413 => "000000000000000000000000",
17414 => "000000000000000000000000",
17415 => "000000000000000000000000",
17416 => "000000000000000000000000",
17417 => "000000000000000000000000",
17418 => "000000000000000000000000",
17419 => "000000000000000000000000",
17420 => "000000000000000000000000",
17421 => "000000000000000000000000",
17422 => "000000000000000000000000",
17423 => "000000000000000000000000",
17424 => "000000000000000000000000",
17425 => "000000000000000000000000",
17426 => "000000000000000000000000",
17427 => "000000000000000000000000",
17428 => "000000000000000000000000",
17429 => "000000000000000000000000",
17430 => "000000000000000000000000",
17431 => "000000000000000000000000",
17432 => "000000000000000000000000",
17433 => "000000000000000000000000",
17434 => "000000000000000000000000",
17435 => "000000000000000000000000",
17436 => "000000000000000000000000",
17437 => "000000000000000000000000",
17438 => "000000000000000000000000",
17439 => "000000000000000000000000",
17440 => "000000000000000000000000",
17441 => "000000000000000000000000",
17442 => "000000000000000000000000",
17443 => "000000000000000000000000",
17444 => "000000000000000000000000",
17445 => "000000000000000000000000",
17446 => "000000000000000000000000",
17447 => "000000000000000000000000",
17448 => "000000000000000000000000",
17449 => "000000000000000000000000",
17450 => "000000000000000000000000",
17451 => "000000000000000000000000",
17452 => "000000000000000000000000",
17453 => "000010100000101000001010",
17454 => "011001100110011001100110",
17455 => "011001100110011001100110",
17456 => "010010100100101001001010",
17457 => "010000110100001101000011",
17458 => "010100010101000101010001",
17459 => "011001100110011001100110",
17460 => "011001000110010001100100",
17461 => "010000110100001101000011",
17462 => "010000110100001101000011",
17463 => "010000110100001101000011",
17464 => "010000110100001101000011",
17465 => "010100000101000001010000",
17466 => "011001100110011001100110",
17467 => "011001010110010101100101",
17468 => "010000110100001101000011",
17469 => "010000110100001101000011",
17470 => "010110110101101101011011",
17471 => "011001100110011001100110",
17472 => "010110100101101001011010",
17473 => "010000110100001101000011",
17474 => "010000110100001101000011",
17475 => "010000110100001101000011",
17476 => "010000110100001101000011",
17477 => "010110100101101001011010",
17478 => "011001100110011001100110",
17479 => "010110110101101101011011",
17480 => "010000110100001101000011",
17481 => "010000110100001101000011",
17482 => "011001100110011001100110",
17483 => "011001100110011001100110",
17484 => "001001100010011000100110",
17485 => "000000000000000000000000",
17486 => "000000000000000000000000",
17487 => "000000000000000000000000",
17488 => "000000000000000000000000",
17489 => "000000000000000000000000",
17490 => "000000000000000000000000",
17491 => "000000000000000000000000",
17492 => "000000000000000000000000",
17493 => "000000000000000000000000",
17494 => "000000000000000000000000",
17495 => "000000000000000000000000",
17496 => "000000000000000000000000",
17497 => "000000000000000000000000",
17498 => "000000000000000000000000",
17499 => "000000000000000000000000",
17500 => "000000000000000000000000",
17501 => "000000000000000000000000",
17502 => "000000000000000000000000",
17503 => "000000000000000000000000",
17504 => "000000000000000000000000",
17505 => "000000000000000000000000",
17506 => "000000000000000000000000",
17507 => "000000000000000000000000",
17508 => "000000000000000000000000",
17509 => "000000000000000000000000",
17510 => "000000000000000000000000",
17511 => "000000000000000000000000",
17512 => "000000000000000000000000",
17513 => "000000000000000000000000",
17514 => "000000000000000000000000",
17515 => "000000000000000000000000",
17516 => "000000000000000000000000",
17517 => "000000000000000000000000",
17518 => "000000000000000000000000",
17519 => "000000000000000000000000",
17520 => "000000000000000000000000",
17521 => "000000000000000000000000",
17522 => "000000000000000000000000",
17523 => "000000000000000000000000",
17524 => "000000000000000000000000",
17525 => "000000000000000000000000",
17526 => "000000000000000000000000",
17527 => "000000000000000000000000",
17528 => "000000000000000000000000",
17529 => "000000000000000000000000",
17530 => "000000000000000000000000",
17531 => "000000000000000000000000",
17532 => "000000000000000000000000",
17533 => "000000000000000000000000",
17534 => "000000000000000000000000",
17535 => "000000000000000000000000",
17536 => "000000000000000000000000",
17537 => "000000000000000000000000",
17538 => "000000000000000000000000",
17539 => "000000000000000000000000",
17540 => "000000000000000000000000",
17541 => "000000000000000000000000",
17542 => "000000000000000000000000",
17543 => "000000000000000000000000",
17544 => "000000000000000000000000",
17545 => "000000000000000000000000",
17546 => "000000000000000000000000",
17547 => "000000000000000000000000",
17548 => "000000000000000000000000",
17549 => "000000000000000000000000",
17550 => "000000000000000000000000",
17551 => "000000000000000000000000",
17552 => "000000000000000000000000",
17553 => "000000000000000000000000",
17554 => "000000000000000000000000",
17555 => "000000000000000000000000",
17556 => "000000000000000000000000",
17557 => "000000000000000000000000",
17558 => "000000000000000000000000",
17559 => "000000000000000000000000",
17560 => "000000000000000000000000",
17561 => "000000000000000000000000",
17562 => "000000000000000000000000",
17563 => "000000000000000000000000",
17564 => "000000000000000000000000",
17565 => "000000000000000000000000",
17566 => "000000000000000000000000",
17567 => "000000000000000000000000",
17568 => "000000000000000000000000",
17569 => "000000000000000000000000",
17570 => "000000000000000000000000",
17571 => "000000000000000000000000",
17572 => "000000000000000000000000",
17573 => "000000000000000000000000",
17574 => "000000000000000000000000",
17575 => "000000000000000000000000",
17576 => "000000000000000000000000",
17577 => "000000000000000000000000",
17578 => "000000000000000000000000",
17579 => "000000000000000000000000",
17580 => "000000000000000000000000",
17581 => "000000000000000000000000",
17582 => "000000000000000000000000",
17583 => "000000000000000000000000",
17584 => "000000000000000000000000",
17585 => "000000000000000000000000",
17586 => "000000000000000000000000",
17587 => "000000000000000000000000",
17588 => "000000000000000000000000",
17589 => "000000000000000000000000",
17590 => "000000000000000000000000",
17591 => "000000000000000000000000",
17592 => "000000000000000000000000",
17593 => "000000000000000000000000",
17594 => "000000000000000000000000",
17595 => "000000000000000000000000",
17596 => "000000000000000000000000",
17597 => "000000000000000000000000",
17598 => "000000000000000000000000",
17599 => "000000000000000000000000",
17600 => "000000000000000000000000",
17601 => "000110100001101000011010",
17602 => "001110110011101100111011",
17603 => "001111000011110000111100",
17604 => "010001110100011101000111",
17605 => "010001110100011101000111",
17606 => "010111000101110001011100",
17607 => "011000100110001001100010",
17608 => "010101110101011101010111",
17609 => "010001110100011101000111",
17610 => "010001110100011101000111",
17611 => "010000110100001101000011",
17612 => "010000110100001101000011",
17613 => "010000110100001101000011",
17614 => "010000110100001101000011",
17615 => "010100000101000001010000",
17616 => "011001100110011001100110",
17617 => "011001010110010101100101",
17618 => "010000110100001101000011",
17619 => "010000110100001101000011",
17620 => "010110110101101101011011",
17621 => "011001100110011001100110",
17622 => "010110100101101001011010",
17623 => "010000110100001101000011",
17624 => "010000110100001101000011",
17625 => "010000110100001101000011",
17626 => "010000110100001101000011",
17627 => "010001100100011001000110",
17628 => "010001110100011101000111",
17629 => "010100000101000001010000",
17630 => "011000100110001001100010",
17631 => "011000100110001001100010",
17632 => "010001110100011101000111",
17633 => "010001110100011101000111",
17634 => "010000000100000001000000",
17635 => "001110110011101100111011",
17636 => "001010100010101000101010",
17637 => "000000000000000000000000",
17638 => "000000000000000000000000",
17639 => "000000000000000000000000",
17640 => "000000000000000000000000",
17641 => "000000000000000000000000",
17642 => "000000000000000000000000",
17643 => "000000000000000000000000",
17644 => "000000000000000000000000",
17645 => "000000000000000000000000",
17646 => "000000000000000000000000",
17647 => "000000000000000000000000",
17648 => "000000000000000000000000",
17649 => "000000000000000000000000",
17650 => "000000000000000000000000",
17651 => "000000000000000000000000",
17652 => "000000000000000000000000",
17653 => "000000000000000000000000",
17654 => "000000000000000000000000",
17655 => "000000000000000000000000",
17656 => "000000000000000000000000",
17657 => "000000000000000000000000",
17658 => "000000000000000000000000",
17659 => "000000000000000000000000",
17660 => "000000000000000000000000",
17661 => "000000000000000000000000",
17662 => "000000000000000000000000",
17663 => "000000000000000000000000",
17664 => "000000000000000000000000",
17665 => "000000000000000000000000",
17666 => "000000000000000000000000",
17667 => "000000000000000000000000",
17668 => "000000000000000000000000",
17669 => "000000000000000000000000",
17670 => "000000000000000000000000",
17671 => "000000000000000000000000",
17672 => "000000000000000000000000",
17673 => "000000000000000000000000",
17674 => "000000000000000000000000",
17675 => "000000000000000000000000",
17676 => "000000000000000000000000",
17677 => "000000000000000000000000",
17678 => "000000000000000000000000",
17679 => "000000000000000000000000",
17680 => "000000000000000000000000",
17681 => "000000000000000000000000",
17682 => "000000000000000000000000",
17683 => "000000000000000000000000",
17684 => "000000000000000000000000",
17685 => "000000000000000000000000",
17686 => "000000000000000000000000",
17687 => "000000000000000000000000",
17688 => "000000000000000000000000",
17689 => "000000000000000000000000",
17690 => "000000000000000000000000",
17691 => "000000000000000000000000",
17692 => "000000000000000000000000",
17693 => "000000000000000000000000",
17694 => "000000000000000000000000",
17695 => "000000000000000000000000",
17696 => "000000000000000000000000",
17697 => "000000000000000000000000",
17698 => "000000000000000000000000",
17699 => "000000000000000000000000",
17700 => "000000000000000000000000",
17701 => "000000000000000000000000",
17702 => "000000000000000000000000",
17703 => "000000000000000000000000",
17704 => "000000000000000000000000",
17705 => "000000000000000000000000",
17706 => "000000000000000000000000",
17707 => "000000000000000000000000",
17708 => "000000000000000000000000",
17709 => "000000000000000000000000",
17710 => "000000000000000000000000",
17711 => "000000000000000000000000",
17712 => "000000000000000000000000",
17713 => "000000000000000000000000",
17714 => "000000000000000000000000",
17715 => "000000000000000000000000",
17716 => "000000000000000000000000",
17717 => "000000000000000000000000",
17718 => "000000000000000000000000",
17719 => "000000000000000000000000",
17720 => "000000000000000000000000",
17721 => "000000000000000000000000",
17722 => "000000000000000000000000",
17723 => "000000000000000000000000",
17724 => "000000000000000000000000",
17725 => "000000000000000000000000",
17726 => "000000000000000000000000",
17727 => "000000000000000000000000",
17728 => "000000000000000000000000",
17729 => "000000000000000000000000",
17730 => "000000000000000000000000",
17731 => "000000000000000000000000",
17732 => "000000000000000000000000",
17733 => "000000000000000000000000",
17734 => "000000000000000000000000",
17735 => "000000000000000000000000",
17736 => "000000000000000000000000",
17737 => "000000000000000000000000",
17738 => "000000000000000000000000",
17739 => "000000000000000000000000",
17740 => "000000000000000000000000",
17741 => "000000000000000000000000",
17742 => "000000000000000000000000",
17743 => "000000000000000000000000",
17744 => "000000000000000000000000",
17745 => "000000000000000000000000",
17746 => "000000000000000000000000",
17747 => "000000000000000000000000",
17748 => "000000000000000000000000",
17749 => "000000000000000000000000",
17750 => "000000000000000000000000",
17751 => "000111010001110100011101",
17752 => "010000110100001101000011",
17753 => "010000110100001101000011",
17754 => "010000110100001101000011",
17755 => "010000110100001101000011",
17756 => "010111110101111101011111",
17757 => "011001100110011001100110",
17758 => "010110000101100001011000",
17759 => "010000110100001101000011",
17760 => "010000110100001101000011",
17761 => "010000110100001101000011",
17762 => "010000110100001101000011",
17763 => "010000110100001101000011",
17764 => "010000110100001101000011",
17765 => "010100000101000001010000",
17766 => "011001100110011001100110",
17767 => "011001010110010101100101",
17768 => "010000110100001101000011",
17769 => "010000110100001101000011",
17770 => "010110110101101101011011",
17771 => "011001100110011001100110",
17772 => "010110100101101001011010",
17773 => "010000110100001101000011",
17774 => "010000110100001101000011",
17775 => "010000110100001101000011",
17776 => "010000110100001101000011",
17777 => "010000110100001101000011",
17778 => "010000110100001101000011",
17779 => "010011100100111001001110",
17780 => "011001100110011001100110",
17781 => "011001100110011001100110",
17782 => "010000110100001101000011",
17783 => "010000110100001101000011",
17784 => "010000110100001101000011",
17785 => "010000110100001101000011",
17786 => "001100000011000000110000",
17787 => "000000000000000000000000",
17788 => "000000000000000000000000",
17789 => "000000000000000000000000",
17790 => "000000000000000000000000",
17791 => "000000000000000000000000",
17792 => "000000000000000000000000",
17793 => "000000000000000000000000",
17794 => "000000000000000000000000",
17795 => "000000000000000000000000",
17796 => "000000000000000000000000",
17797 => "000000000000000000000000",
17798 => "000000000000000000000000",
17799 => "000000000000000000000000",
17800 => "000000000000000000000000",
17801 => "000000000000000000000000",
17802 => "000000000000000000000000",
17803 => "000000000000000000000000",
17804 => "000000000000000000000000",
17805 => "000000000000000000000000",
17806 => "000000000000000000000000",
17807 => "000000000000000000000000",
17808 => "000000000000000000000000",
17809 => "000000000000000000000000",
17810 => "000000000000000000000000",
17811 => "000000000000000000000000",
17812 => "000000000000000000000000",
17813 => "000000000000000000000000",
17814 => "000000000000000000000000",
17815 => "000000000000000000000000",
17816 => "000000000000000000000000",
17817 => "000000000000000000000000",
17818 => "000000000000000000000000",
17819 => "000000000000000000000000",
17820 => "000000000000000000000000",
17821 => "000000000000000000000000",
17822 => "000000000000000000000000",
17823 => "000000000000000000000000",
17824 => "000000000000000000000000",
17825 => "000000000000000000000000",
17826 => "000000000000000000000000",
17827 => "000000000000000000000000",
17828 => "000000000000000000000000",
17829 => "000000000000000000000000",
17830 => "000000000000000000000000",
17831 => "000000000000000000000000",
17832 => "000000000000000000000000",
17833 => "000000000000000000000000",
17834 => "000000000000000000000000",
17835 => "000000000000000000000000",
17836 => "000000000000000000000000",
17837 => "000000000000000000000000",
17838 => "000000000000000000000000",
17839 => "000000000000000000000000",
17840 => "000000000000000000000000",
17841 => "000000000000000000000000",
17842 => "000000000000000000000000",
17843 => "000000000000000000000000",
17844 => "000000000000000000000000",
17845 => "000000000000000000000000",
17846 => "000000000000000000000000",
17847 => "000000000000000000000000",
17848 => "000000000000000000000000",
17849 => "000000000000000000000000",
17850 => "000000000000000000000000",
17851 => "000000000000000000000000",
17852 => "000000000000000000000000",
17853 => "000000000000000000000000",
17854 => "000000000000000000000000",
17855 => "000000000000000000000000",
17856 => "000000000000000000000000",
17857 => "000000000000000000000000",
17858 => "000000000000000000000000",
17859 => "000000000000000000000000",
17860 => "000000000000000000000000",
17861 => "000000000000000000000000",
17862 => "000000000000000000000000",
17863 => "000000000000000000000000",
17864 => "000000000000000000000000",
17865 => "000000000000000000000000",
17866 => "000000000000000000000000",
17867 => "000000000000000000000000",
17868 => "000000000000000000000000",
17869 => "000000000000000000000000",
17870 => "000000000000000000000000",
17871 => "000000000000000000000000",
17872 => "000000000000000000000000",
17873 => "000000000000000000000000",
17874 => "000000000000000000000000",
17875 => "000000000000000000000000",
17876 => "000000000000000000000000",
17877 => "000000000000000000000000",
17878 => "000000000000000000000000",
17879 => "000000000000000000000000",
17880 => "000000000000000000000000",
17881 => "000000000000000000000000",
17882 => "000000000000000000000000",
17883 => "000000000000000000000000",
17884 => "000000000000000000000000",
17885 => "000000000000000000000000",
17886 => "000000000000000000000000",
17887 => "000000000000000000000000",
17888 => "000000000000000000000000",
17889 => "000000000000000000000000",
17890 => "000000000000000000000000",
17891 => "000000000000000000000000",
17892 => "000000000000000000000000",
17893 => "000000000000000000000000",
17894 => "000000000000000000000000",
17895 => "000000000000000000000000",
17896 => "000000000000000000000000",
17897 => "000000000000000000000000",
17898 => "000000000000000000000000",
17899 => "000110100001101000011010",
17900 => "000111110001111100011111",
17901 => "001011110010111100101111",
17902 => "010000110100001101000011",
17903 => "010000110100001101000011",
17904 => "010000110100001101000011",
17905 => "010000110100001101000011",
17906 => "010111110101111101011111",
17907 => "011001100110011001100110",
17908 => "010010110100101101001011",
17909 => "001001000010010000100100",
17910 => "001001000010010000100100",
17911 => "001001000010010000100100",
17912 => "001001000010010000100100",
17913 => "001001000010010000100100",
17914 => "001001000010010000100100",
17915 => "001111000011110000111100",
17916 => "011001100110011001100110",
17917 => "011001010110010101100101",
17918 => "010100110101001101010011",
17919 => "010100110101001101010011",
17920 => "001111110011111100111111",
17921 => "001101100011011000110110",
17922 => "001100000011000000110000",
17923 => "001001000010010000100100",
17924 => "001001000010010000100100",
17925 => "001001000010010000100100",
17926 => "001001000010010000100100",
17927 => "001001000010010000100100",
17928 => "001001000010010000100100",
17929 => "001110000011100000111000",
17930 => "011001100110011001100110",
17931 => "011001100110011001100110",
17932 => "010000110100001101000011",
17933 => "010000110100001101000011",
17934 => "010000110100001101000011",
17935 => "010000110100001101000011",
17936 => "001110010011100100111001",
17937 => "000111110001111100011111",
17938 => "000111110001111100011111",
17939 => "000000000000000000000000",
17940 => "000000000000000000000000",
17941 => "000000000000000000000000",
17942 => "000000000000000000000000",
17943 => "000000000000000000000000",
17944 => "000000000000000000000000",
17945 => "000000000000000000000000",
17946 => "000000000000000000000000",
17947 => "000000000000000000000000",
17948 => "000000000000000000000000",
17949 => "000000000000000000000000",
17950 => "000000000000000000000000",
17951 => "000000000000000000000000",
17952 => "000000000000000000000000",
17953 => "000000000000000000000000",
17954 => "000000000000000000000000",
17955 => "000000000000000000000000",
17956 => "000000000000000000000000",
17957 => "000000000000000000000000",
17958 => "000000000000000000000000",
17959 => "000000000000000000000000",
17960 => "000000000000000000000000",
17961 => "000000000000000000000000",
17962 => "000000000000000000000000",
17963 => "000000000000000000000000",
17964 => "000000000000000000000000",
17965 => "000000000000000000000000",
17966 => "000000000000000000000000",
17967 => "000000000000000000000000",
17968 => "000000000000000000000000",
17969 => "000000000000000000000000",
17970 => "000000000000000000000000",
17971 => "000000000000000000000000",
17972 => "000000000000000000000000",
17973 => "000000000000000000000000",
17974 => "000000000000000000000000",
17975 => "000000000000000000000000",
17976 => "000000000000000000000000",
17977 => "000000000000000000000000",
17978 => "000000000000000000000000",
17979 => "000000000000000000000000",
17980 => "000000000000000000000000",
17981 => "000000000000000000000000",
17982 => "000000000000000000000000",
17983 => "000000000000000000000000",
17984 => "000000000000000000000000",
17985 => "000000000000000000000000",
17986 => "000000000000000000000000",
17987 => "000000000000000000000000",
17988 => "000000000000000000000000",
17989 => "000000000000000000000000",
17990 => "000000000000000000000000",
17991 => "000000000000000000000000",
17992 => "000000000000000000000000",
17993 => "000000000000000000000000",
17994 => "000000000000000000000000",
17995 => "000000000000000000000000",
17996 => "000000000000000000000000",
17997 => "000000000000000000000000",
17998 => "000000000000000000000000",
17999 => "000000000000000000000000",
18000 => "000000000000000000000000",
18001 => "000000000000000000000000",
18002 => "000000000000000000000000",
18003 => "000000000000000000000000",
18004 => "000000000000000000000000",
18005 => "000000000000000000000000",
18006 => "000000000000000000000000",
18007 => "000000000000000000000000",
18008 => "000000000000000000000000",
18009 => "000000000000000000000000",
18010 => "000000000000000000000000",
18011 => "000000000000000000000000",
18012 => "000000000000000000000000",
18013 => "000000000000000000000000",
18014 => "000000000000000000000000",
18015 => "000000000000000000000000",
18016 => "000000000000000000000000",
18017 => "000000000000000000000000",
18018 => "000000000000000000000000",
18019 => "000000000000000000000000",
18020 => "000000000000000000000000",
18021 => "000000000000000000000000",
18022 => "000000000000000000000000",
18023 => "000000000000000000000000",
18024 => "000000000000000000000000",
18025 => "000000000000000000000000",
18026 => "000000000000000000000000",
18027 => "000000000000000000000000",
18028 => "000000000000000000000000",
18029 => "000000000000000000000000",
18030 => "000000000000000000000000",
18031 => "000000000000000000000000",
18032 => "000000000000000000000000",
18033 => "000000000000000000000000",
18034 => "000000000000000000000000",
18035 => "000000000000000000000000",
18036 => "000000000000000000000000",
18037 => "000000000000000000000000",
18038 => "000000000000000000000000",
18039 => "000000000000000000000000",
18040 => "000000000000000000000000",
18041 => "000000000000000000000000",
18042 => "000000000000000000000000",
18043 => "000000000000000000000000",
18044 => "000000000000000000000000",
18045 => "000000000000000000000000",
18046 => "000000000000000000000000",
18047 => "000000000000000000000000",
18048 => "000000000000000000000000",
18049 => "001110000011100000111000",
18050 => "010000110100001101000011",
18051 => "010000110100001101000011",
18052 => "010000110100001101000011",
18053 => "010000110100001101000011",
18054 => "010000110100001101000011",
18055 => "010000110100001101000011",
18056 => "010111110101111101011111",
18057 => "011001100110011001100110",
18058 => "001111010011110100111101",
18059 => "000000000000000000000000",
18060 => "000000000000000000000000",
18061 => "000000000000000000000000",
18062 => "000000000000000000000000",
18063 => "000000000000000000000000",
18064 => "000000000000000000000000",
18065 => "001001100010011000100110",
18066 => "011001100110011001100110",
18067 => "011001100110011001100110",
18068 => "011001100110011001100110",
18069 => "011001100110011001100110",
18070 => "001000000010000000100000",
18071 => "000000000000000000000000",
18072 => "000000000000000000000000",
18073 => "000000000000000000000000",
18074 => "000000000000000000000000",
18075 => "000000000000000000000000",
18076 => "000000000000000000000000",
18077 => "000000000000000000000000",
18078 => "000000000000000000000000",
18079 => "001000000010000000100000",
18080 => "011001100110011001100110",
18081 => "011001100110011001100110",
18082 => "010000110100001101000011",
18083 => "010000110100001101000011",
18084 => "010000110100001101000011",
18085 => "010000110100001101000011",
18086 => "010000110100001101000011",
18087 => "010000110100001101000011",
18088 => "010000110100001101000011",
18089 => "000000010000000100000001",
18090 => "000000000000000000000000",
18091 => "000000000000000000000000",
18092 => "000000000000000000000000",
18093 => "000000000000000000000000",
18094 => "000000000000000000000000",
18095 => "000000000000000000000000",
18096 => "000000000000000000000000",
18097 => "000000000000000000000000",
18098 => "000000000000000000000000",
18099 => "000000000000000000000000",
18100 => "000000000000000000000000",
18101 => "000000000000000000000000",
18102 => "000000000000000000000000",
18103 => "000000000000000000000000",
18104 => "000000000000000000000000",
18105 => "000000000000000000000000",
18106 => "000000000000000000000000",
18107 => "000000000000000000000000",
18108 => "000000000000000000000000",
18109 => "000000000000000000000000",
18110 => "000000000000000000000000",
18111 => "000000000000000000000000",
18112 => "000000000000000000000000",
18113 => "000000000000000000000000",
18114 => "000000000000000000000000",
18115 => "000000000000000000000000",
18116 => "000000000000000000000000",
18117 => "000000000000000000000000",
18118 => "000000000000000000000000",
18119 => "000000000000000000000000",
18120 => "000000000000000000000000",
18121 => "000000000000000000000000",
18122 => "000000000000000000000000",
18123 => "000000000000000000000000",
18124 => "000000000000000000000000",
18125 => "000000000000000000000000",
18126 => "000000000000000000000000",
18127 => "000000000000000000000000",
18128 => "000000000000000000000000",
18129 => "000000000000000000000000",
18130 => "000000000000000000000000",
18131 => "000000000000000000000000",
18132 => "000000000000000000000000",
18133 => "000000000000000000000000",
18134 => "000000000000000000000000",
18135 => "000000000000000000000000",
18136 => "000000000000000000000000",
18137 => "000000000000000000000000",
18138 => "000000000000000000000000",
18139 => "000000000000000000000000",
18140 => "000000000000000000000000",
18141 => "000000000000000000000000",
18142 => "000000000000000000000000",
18143 => "000000000000000000000000",
18144 => "000000000000000000000000",
18145 => "000000000000000000000000",
18146 => "000000000000000000000000",
18147 => "000000000000000000000000",
18148 => "000000000000000000000000",
18149 => "000000000000000000000000",
18150 => "000000000000000000000000",
18151 => "000000000000000000000000",
18152 => "000000000000000000000000",
18153 => "000000000000000000000000",
18154 => "000000000000000000000000",
18155 => "000000000000000000000000",
18156 => "000000000000000000000000",
18157 => "000000000000000000000000",
18158 => "000000000000000000000000",
18159 => "000000000000000000000000",
18160 => "000000000000000000000000",
18161 => "000000000000000000000000",
18162 => "000000000000000000000000",
18163 => "000000000000000000000000",
18164 => "000000000000000000000000",
18165 => "000000000000000000000000",
18166 => "000000000000000000000000",
18167 => "000000000000000000000000",
18168 => "000000000000000000000000",
18169 => "000000000000000000000000",
18170 => "000000000000000000000000",
18171 => "000000000000000000000000",
18172 => "000000000000000000000000",
18173 => "000000000000000000000000",
18174 => "000000000000000000000000",
18175 => "000000000000000000000000",
18176 => "000000000000000000000000",
18177 => "000000000000000000000000",
18178 => "000000000000000000000000",
18179 => "000000000000000000000000",
18180 => "000000000000000000000000",
18181 => "000000000000000000000000",
18182 => "000000000000000000000000",
18183 => "000000000000000000000000",
18184 => "000000000000000000000000",
18185 => "000000000000000000000000",
18186 => "000000000000000000000000",
18187 => "000000000000000000000000",
18188 => "000000000000000000000000",
18189 => "000000000000000000000000",
18190 => "000000000000000000000000",
18191 => "000000000000000000000000",
18192 => "000000000000000000000000",
18193 => "000000000000000000000000",
18194 => "000000000000000000000000",
18195 => "000000000000000000000000",
18196 => "000000010000000100000001",
18197 => "000010000000100000001000",
18198 => "000010000000100000001000",
18199 => "001110010011100100111001",
18200 => "010000110100001101000011",
18201 => "010000110100001101000011",
18202 => "010000110100001101000011",
18203 => "010000110100001101000011",
18204 => "010000110100001101000011",
18205 => "010000110100001101000011",
18206 => "010101010101010101010101",
18207 => "010110010101100101011001",
18208 => "001110110011101000110101",
18209 => "000100000000110000000000",
18210 => "000100000000110000000001",
18211 => "000011010000110100001101",
18212 => "000011010000110100001101",
18213 => "000011110000110000000011",
18214 => "000100000000110000000000",
18215 => "001100000010111000100110",
18216 => "011001100110011001100110",
18217 => "011001100110011001100110",
18218 => "010110010101100101011001",
18219 => "010110010101100101011001",
18220 => "001001010010010100100101",
18221 => "000011010000110100001101",
18222 => "000011100000110000001000",
18223 => "000100000000110000000000",
18224 => "000100000000110000000000",
18225 => "000011010000110100001101",
18226 => "000011010000110100001101",
18227 => "000011110000110000000100",
18228 => "000100000000110000000000",
18229 => "001001110010010000011100",
18230 => "010110010101100101011001",
18231 => "010110010101100101011001",
18232 => "010000110100001101000011",
18233 => "010000110100001101000011",
18234 => "010000110100001101000011",
18235 => "010000110100001101000011",
18236 => "010000110100001101000011",
18237 => "010000110100001101000011",
18238 => "010000110100001101000011",
18239 => "000010010000100100001001",
18240 => "000010000000100000001000",
18241 => "000000110000001100000011",
18242 => "000000000000000000000000",
18243 => "000000000000000000000000",
18244 => "000000000000000000000000",
18245 => "000000000000000000000000",
18246 => "000000000000000000000000",
18247 => "000000000000000000000000",
18248 => "000000000000000000000000",
18249 => "000000000000000000000000",
18250 => "000000000000000000000000",
18251 => "000000000000000000000000",
18252 => "000000000000000000000000",
18253 => "000000000000000000000000",
18254 => "000000000000000000000000",
18255 => "000000000000000000000000",
18256 => "000000000000000000000000",
18257 => "000000000000000000000000",
18258 => "000000000000000000000000",
18259 => "000000000000000000000000",
18260 => "000000000000000000000000",
18261 => "000000000000000000000000",
18262 => "000000000000000000000000",
18263 => "000000000000000000000000",
18264 => "000000000000000000000000",
18265 => "000000000000000000000000",
18266 => "000000000000000000000000",
18267 => "000000000000000000000000",
18268 => "000000000000000000000000",
18269 => "000000000000000000000000",
18270 => "000000000000000000000000",
18271 => "000000000000000000000000",
18272 => "000000000000000000000000",
18273 => "000000000000000000000000",
18274 => "000000000000000000000000",
18275 => "000000000000000000000000",
18276 => "000000000000000000000000",
18277 => "000000000000000000000000",
18278 => "000000000000000000000000",
18279 => "000000000000000000000000",
18280 => "000000000000000000000000",
18281 => "000000000000000000000000",
18282 => "000000000000000000000000",
18283 => "000000000000000000000000",
18284 => "000000000000000000000000",
18285 => "000000000000000000000000",
18286 => "000000000000000000000000",
18287 => "000000000000000000000000",
18288 => "000000000000000000000000",
18289 => "000000000000000000000000",
18290 => "000000000000000000000000",
18291 => "000000000000000000000000",
18292 => "000000000000000000000000",
18293 => "000000000000000000000000",
18294 => "000000000000000000000000",
18295 => "000000000000000000000000",
18296 => "000000000000000000000000",
18297 => "000000000000000000000000",
18298 => "000000000000000000000000",
18299 => "000000000000000000000000",
18300 => "000000000000000000000000",
18301 => "000000000000000000000000",
18302 => "000000000000000000000000",
18303 => "000000000000000000000000",
18304 => "000000000000000000000000",
18305 => "000000000000000000000000",
18306 => "000000000000000000000000",
18307 => "000000000000000000000000",
18308 => "000000000000000000000000",
18309 => "000000000000000000000000",
18310 => "000000000000000000000000",
18311 => "000000000000000000000000",
18312 => "000000000000000000000000",
18313 => "000000000000000000000000",
18314 => "000000000000000000000000",
18315 => "000000000000000000000000",
18316 => "000000000000000000000000",
18317 => "000000000000000000000000",
18318 => "000000000000000000000000",
18319 => "000000000000000000000000",
18320 => "000000000000000000000000",
18321 => "000000000000000000000000",
18322 => "000000000000000000000000",
18323 => "000000000000000000000000",
18324 => "000000000000000000000000",
18325 => "000000000000000000000000",
18326 => "000000000000000000000000",
18327 => "000000000000000000000000",
18328 => "000000000000000000000000",
18329 => "000000000000000000000000",
18330 => "000000000000000000000000",
18331 => "000000000000000000000000",
18332 => "000000000000000000000000",
18333 => "000000000000000000000000",
18334 => "000000000000000000000000",
18335 => "000000000000000000000000",
18336 => "000000000000000000000000",
18337 => "000000000000000000000000",
18338 => "000000000000000000000000",
18339 => "000000000000000000000000",
18340 => "000000000000000000000000",
18341 => "000000000000000000000000",
18342 => "000000000000000000000000",
18343 => "000000000000000000000000",
18344 => "000000000000000000000000",
18345 => "000000000000000000000000",
18346 => "000010000000100000001000",
18347 => "010000110100001101000011",
18348 => "010000110100001101000011",
18349 => "010000110100001101000011",
18350 => "010000110100001101000011",
18351 => "010000110100001101000011",
18352 => "010000110100001101000011",
18353 => "010000110100001101000011",
18354 => "010000110100001101000011",
18355 => "010000110100001101000011",
18356 => "000011100000111000001110",
18357 => "000000000000000000000000",
18358 => "001101000010011100000000",
18359 => "011111110110000000000000",
18360 => "011111010110000000000110",
18361 => "011001100110011001100110",
18362 => "011001100110011001100110",
18363 => "011110000110001000011100",
18364 => "011111110110000000000000",
18365 => "011101100110001000100110",
18366 => "011001100110011001100110",
18367 => "011000110110001101100011",
18368 => "000000000000000000000000",
18369 => "000000000000000000000000",
18370 => "010001100100011001000110",
18371 => "011001100110011001100110",
18372 => "011011110110010001000011",
18373 => "011111110110000000000000",
18374 => "011111110110000000000000",
18375 => "011001100110011001100110",
18376 => "011001100110011001100110",
18377 => "011101100110001000100011",
18378 => "011111110110000000000000",
18379 => "010101110100001000000000",
18380 => "000000000000000000000000",
18381 => "000000000000000000000000",
18382 => "010000110100001101000011",
18383 => "010000110100001101000011",
18384 => "010000110100001101000011",
18385 => "010000110100001101000011",
18386 => "010000110100001101000011",
18387 => "010000110100001101000011",
18388 => "010000110100001101000011",
18389 => "010000110100001101000011",
18390 => "010000110100001101000011",
18391 => "000110110001101100011011",
18392 => "000000000000000000000000",
18393 => "000000000000000000000000",
18394 => "000000000000000000000000",
18395 => "000000000000000000000000",
18396 => "000000000000000000000000",
18397 => "000000000000000000000000",
18398 => "000000000000000000000000",
18399 => "000000000000000000000000",
18400 => "000000000000000000000000",
18401 => "000000000000000000000000",
18402 => "000000000000000000000000",
18403 => "000000000000000000000000",
18404 => "000000000000000000000000",
18405 => "000000000000000000000000",
18406 => "000000000000000000000000",
18407 => "000000000000000000000000",
18408 => "000000000000000000000000",
18409 => "000000000000000000000000",
18410 => "000000000000000000000000",
18411 => "000000000000000000000000",
18412 => "000000000000000000000000",
18413 => "000000000000000000000000",
18414 => "000000000000000000000000",
18415 => "000000000000000000000000",
18416 => "000000000000000000000000",
18417 => "000000000000000000000000",
18418 => "000000000000000000000000",
18419 => "000000000000000000000000",
18420 => "000000000000000000000000",
18421 => "000000000000000000000000",
18422 => "000000000000000000000000",
18423 => "000000000000000000000000",
18424 => "000000000000000000000000",
18425 => "000000000000000000000000",
18426 => "000000000000000000000000",
18427 => "000000000000000000000000",
18428 => "000000000000000000000000",
18429 => "000000000000000000000000",
18430 => "000000000000000000000000",
18431 => "000000000000000000000000",
18432 => "000000000000000000000000",
18433 => "000000000000000000000000",
18434 => "000000000000000000000000",
18435 => "000000000000000000000000",
18436 => "000000000000000000000000",
18437 => "000000000000000000000000",
18438 => "000000000000000000000000",
18439 => "000000000000000000000000",
18440 => "000000000000000000000000",
18441 => "000000000000000000000000",
18442 => "000000000000000000000000",
18443 => "000000000000000000000000",
18444 => "000000000000000000000000",
18445 => "000000000000000000000000",
18446 => "000000000000000000000000",
18447 => "000000000000000000000000",
18448 => "000000000000000000000000",
18449 => "000000000000000000000000",
18450 => "000000000000000000000000",
18451 => "000000000000000000000000",
18452 => "000000000000000000000000",
18453 => "000000000000000000000000",
18454 => "000000000000000000000000",
18455 => "000000000000000000000000",
18456 => "000000000000000000000000",
18457 => "000000000000000000000000",
18458 => "000000000000000000000000",
18459 => "000000000000000000000000",
18460 => "000000000000000000000000",
18461 => "000000000000000000000000",
18462 => "000000000000000000000000",
18463 => "000000000000000000000000",
18464 => "000000000000000000000000",
18465 => "000000000000000000000000",
18466 => "000000000000000000000000",
18467 => "000000000000000000000000",
18468 => "000000000000000000000000",
18469 => "000000000000000000000000",
18470 => "000000000000000000000000",
18471 => "000000000000000000000000",
18472 => "000000000000000000000000",
18473 => "000000000000000000000000",
18474 => "000000000000000000000000",
18475 => "000000000000000000000000",
18476 => "000000000000000000000000",
18477 => "000000000000000000000000",
18478 => "000000000000000000000000",
18479 => "000000000000000000000000",
18480 => "000000000000000000000000",
18481 => "000000000000000000000000",
18482 => "000000000000000000000000",
18483 => "000000000000000000000000",
18484 => "000000000000000000000000",
18485 => "000000000000000000000000",
18486 => "000000000000000000000000",
18487 => "000000000000000000000000",
18488 => "000000000000000000000000",
18489 => "000000000000000000000000",
18490 => "000000000000000000000000",
18491 => "000000000000000000000000",
18492 => "000000000000000000000000",
18493 => "000000000000000000000000",
18494 => "000000000000000000000000",
18495 => "000000000000000000000000",
18496 => "000010000000100000001000",
18497 => "010000110100001101000011",
18498 => "010000110100001101000011",
18499 => "010000110100001101000011",
18500 => "010000110100001101000011",
18501 => "010000110100001101000011",
18502 => "010000110100001101000011",
18503 => "010000110100001101000011",
18504 => "010000110100001101000011",
18505 => "010000110100001101000011",
18506 => "000011100000111000001110",
18507 => "000000000000000000000000",
18508 => "001101000010011100000000",
18509 => "011111110110000000000000",
18510 => "011111010110000000000110",
18511 => "011001100110011001100110",
18512 => "011001100110011001100110",
18513 => "011110000110001000011100",
18514 => "011111110110000000000000",
18515 => "011101100110001000100110",
18516 => "011001100110011001100110",
18517 => "011000110110001101100011",
18518 => "000000000000000000000000",
18519 => "000000000000000000000000",
18520 => "010001100100011001000110",
18521 => "011001100110011001100110",
18522 => "011011110110010001000011",
18523 => "011111110110000000000000",
18524 => "011111110110000000000000",
18525 => "011001100110011001100110",
18526 => "011001100110011001100110",
18527 => "011101100110001000100011",
18528 => "011111110110000000000000",
18529 => "010101110100001000000000",
18530 => "000000000000000000000000",
18531 => "000000000000000000000000",
18532 => "010000110100001101000011",
18533 => "010000110100001101000011",
18534 => "010000110100001101000011",
18535 => "010000110100001101000011",
18536 => "010000110100001101000011",
18537 => "010000110100001101000011",
18538 => "010000110100001101000011",
18539 => "010000110100001101000011",
18540 => "010000110100001101000011",
18541 => "000110110001101100011011",
18542 => "000000000000000000000000",
18543 => "000000000000000000000000",
18544 => "000000000000000000000000",
18545 => "000000000000000000000000",
18546 => "000000000000000000000000",
18547 => "000000000000000000000000",
18548 => "000000000000000000000000",
18549 => "000000000000000000000000",
18550 => "000000000000000000000000",
18551 => "000000000000000000000000",
18552 => "000000000000000000000000",
18553 => "000000000000000000000000",
18554 => "000000000000000000000000",
18555 => "000000000000000000000000",
18556 => "000000000000000000000000",
18557 => "000000000000000000000000",
18558 => "000000000000000000000000",
18559 => "000000000000000000000000",
18560 => "000000000000000000000000",
18561 => "000000000000000000000000",
18562 => "000000000000000000000000",
18563 => "000000000000000000000000",
18564 => "000000000000000000000000",
18565 => "000000000000000000000000",
18566 => "000000000000000000000000",
18567 => "000000000000000000000000",
18568 => "000000000000000000000000",
18569 => "000000000000000000000000",
18570 => "000000000000000000000000",
18571 => "000000000000000000000000",
18572 => "000000000000000000000000",
18573 => "000000000000000000000000",
18574 => "000000000000000000000000",
18575 => "000000000000000000000000",
18576 => "000000000000000000000000",
18577 => "000000000000000000000000",
18578 => "000000000000000000000000",
18579 => "000000000000000000000000",
18580 => "000000000000000000000000",
18581 => "000000000000000000000000",
18582 => "000000000000000000000000",
18583 => "000000000000000000000000",
18584 => "000000000000000000000000",
18585 => "000000000000000000000000",
18586 => "000000000000000000000000",
18587 => "000000000000000000000000",
18588 => "000000000000000000000000",
18589 => "000000000000000000000000",
18590 => "000000000000000000000000",
18591 => "000000000000000000000000",
18592 => "000000000000000000000000",
18593 => "000000000000000000000000",
18594 => "000000000000000000000000",
18595 => "000000000000000000000000",
18596 => "000000000000000000000000",
18597 => "000000000000000000000000",
18598 => "000000000000000000000000",
18599 => "000000000000000000000000",
18600 => "000000000000000000000000",
18601 => "000000000000000000000000",
18602 => "000000000000000000000000",
18603 => "000000000000000000000000",
18604 => "000000000000000000000000",
18605 => "000000000000000000000000",
18606 => "000000000000000000000000",
18607 => "000000000000000000000000",
18608 => "000000000000000000000000",
18609 => "000000000000000000000000",
18610 => "000000000000000000000000",
18611 => "000000000000000000000000",
18612 => "000000000000000000000000",
18613 => "000000000000000000000000",
18614 => "000000000000000000000000",
18615 => "000000000000000000000000",
18616 => "000000000000000000000000",
18617 => "000000000000000000000000",
18618 => "000000000000000000000000",
18619 => "000000000000000000000000",
18620 => "000000000000000000000000",
18621 => "000000000000000000000000",
18622 => "000000000000000000000000",
18623 => "000000000000000000000000",
18624 => "000000000000000000000000",
18625 => "000000000000000000000000",
18626 => "000000000000000000000000",
18627 => "000000000000000000000000",
18628 => "000000000000000000000000",
18629 => "000000000000000000000000",
18630 => "000000000000000000000000",
18631 => "000000000000000000000000",
18632 => "000000000000000000000000",
18633 => "000000000000000000000000",
18634 => "000000000000000000000000",
18635 => "000000000000000000000000",
18636 => "000000000000000000000000",
18637 => "000000000000000000000000",
18638 => "000000000000000000000000",
18639 => "000000000000000000000000",
18640 => "000000000000000000000000",
18641 => "000000000000000000000000",
18642 => "000000000000000000000000",
18643 => "000000000000000000000000",
18644 => "000110100001101000011010",
18645 => "001110000011100000111000",
18646 => "001110010011100100111001",
18647 => "010000110100001101000011",
18648 => "010000110100001101000011",
18649 => "010000110100001101000011",
18650 => "010000110100001101000011",
18651 => "010000110100001101000011",
18652 => "010000110100001101000011",
18653 => "010000110100001101000011",
18654 => "010000110100001101000011",
18655 => "010000110100001101000011",
18656 => "000011100000111000001110",
18657 => "000000000000000000000000",
18658 => "001101000010011100000000",
18659 => "011111110110000000000000",
18660 => "011111010110000000000110",
18661 => "011001100110011001100110",
18662 => "011001100110011001100110",
18663 => "011110000110001000011100",
18664 => "011111110110000000000000",
18665 => "011101100110001000100110",
18666 => "011001100110011001100110",
18667 => "011000110110001101100011",
18668 => "000000000000000000000000",
18669 => "000000000000000000000000",
18670 => "010001100100011001000110",
18671 => "011001100110011001100110",
18672 => "011011110110010001000011",
18673 => "011111110110000000000000",
18674 => "011111110110000000000000",
18675 => "011001100110011001100110",
18676 => "011001100110011001100110",
18677 => "011101100110001000100011",
18678 => "011111110110000000000000",
18679 => "010101110100001000000000",
18680 => "000000000000000000000000",
18681 => "000000000000000000000000",
18682 => "010000110100001101000011",
18683 => "010000110100001101000011",
18684 => "010000110100001101000011",
18685 => "010000110100001101000011",
18686 => "010000110100001101000011",
18687 => "010000110100001101000011",
18688 => "010000110100001101000011",
18689 => "010000110100001101000011",
18690 => "010000110100001101000011",
18691 => "001111010011110100111101",
18692 => "001110000011100000111000",
18693 => "001010100010101000101010",
18694 => "000000000000000000000000",
18695 => "000000000000000000000000",
18696 => "000000000000000000000000",
18697 => "000000000000000000000000",
18698 => "000000000000000000000000",
18699 => "000000000000000000000000",
18700 => "000000000000000000000000",
18701 => "000000000000000000000000",
18702 => "000000000000000000000000",
18703 => "000000000000000000000000",
18704 => "000000000000000000000000",
18705 => "000000000000000000000000",
18706 => "000000000000000000000000",
18707 => "000000000000000000000000",
18708 => "000000000000000000000000",
18709 => "000000000000000000000000",
18710 => "000000000000000000000000",
18711 => "000000000000000000000000",
18712 => "000000000000000000000000",
18713 => "000000000000000000000000",
18714 => "000000000000000000000000",
18715 => "000000000000000000000000",
18716 => "000000000000000000000000",
18717 => "000000000000000000000000",
18718 => "000000000000000000000000",
18719 => "000000000000000000000000",
18720 => "000000000000000000000000",
18721 => "000000000000000000000000",
18722 => "000000000000000000000000",
18723 => "000000000000000000000000",
18724 => "000000000000000000000000",
18725 => "000000000000000000000000",
18726 => "000000000000000000000000",
18727 => "000000000000000000000000",
18728 => "000000000000000000000000",
18729 => "000000000000000000000000",
18730 => "000000000000000000000000",
18731 => "000000000000000000000000",
18732 => "000000000000000000000000",
18733 => "000000000000000000000000",
18734 => "000000000000000000000000",
18735 => "000000000000000000000000",
18736 => "000000000000000000000000",
18737 => "000000000000000000000000",
18738 => "000000000000000000000000",
18739 => "000000000000000000000000",
18740 => "000000000000000000000000",
18741 => "000000000000000000000000",
18742 => "000000000000000000000000",
18743 => "000000000000000000000000",
18744 => "000000000000000000000000",
18745 => "000000000000000000000000",
18746 => "000000000000000000000000",
18747 => "000000000000000000000000",
18748 => "000000000000000000000000",
18749 => "000000000000000000000000",
18750 => "000000000000000000000000",
18751 => "000000000000000000000000",
18752 => "000000000000000000000000",
18753 => "000000000000000000000000",
18754 => "000000000000000000000000",
18755 => "000000000000000000000000",
18756 => "000000000000000000000000",
18757 => "000000000000000000000000",
18758 => "000000000000000000000000",
18759 => "000000000000000000000000",
18760 => "000000000000000000000000",
18761 => "000000000000000000000000",
18762 => "000000000000000000000000",
18763 => "000000000000000000000000",
18764 => "000000000000000000000000",
18765 => "000000000000000000000000",
18766 => "000000000000000000000000",
18767 => "000000000000000000000000",
18768 => "000000000000000000000000",
18769 => "000000000000000000000000",
18770 => "000000000000000000000000",
18771 => "000000000000000000000000",
18772 => "000000000000000000000000",
18773 => "000000000000000000000000",
18774 => "000000000000000000000000",
18775 => "000000000000000000000000",
18776 => "000000000000000000000000",
18777 => "000000000000000000000000",
18778 => "000000000000000000000000",
18779 => "000000000000000000000000",
18780 => "000000000000000000000000",
18781 => "000000000000000000000000",
18782 => "000000000000000000000000",
18783 => "000000000000000000000000",
18784 => "000000000000000000000000",
18785 => "000000000000000000000000",
18786 => "000000000000000000000000",
18787 => "000000000000000000000000",
18788 => "000000000000000000000000",
18789 => "000000000000000000000000",
18790 => "000000000000000000000000",
18791 => "000000000000000000000000",
18792 => "000000000000000000000000",
18793 => "000000000000000000000000",
18794 => "000111110001111100011111",
18795 => "010000110100001101000011",
18796 => "010000110100001101000011",
18797 => "010000110100001101000011",
18798 => "010000110100001101000011",
18799 => "010000110100001101000011",
18800 => "010000110100001101000011",
18801 => "010000110100001101000011",
18802 => "010000110100001101000011",
18803 => "010000110100001101000011",
18804 => "010000110100001101000011",
18805 => "010000110100001101000011",
18806 => "000011100000111000001110",
18807 => "000000000000000000000000",
18808 => "001101000010011100000000",
18809 => "011111110110000000000000",
18810 => "011111010110000000000110",
18811 => "011001100110011001100110",
18812 => "011001100110011001100110",
18813 => "011110000110001000011100",
18814 => "011111110110000000000000",
18815 => "011101100110001000100110",
18816 => "011001100110011001100110",
18817 => "011000110110001101100011",
18818 => "000000000000000000000000",
18819 => "000000000000000000000000",
18820 => "010001100100011001000110",
18821 => "011001100110011001100110",
18822 => "011011110110010001000011",
18823 => "011111110110000000000000",
18824 => "011111110110000000000000",
18825 => "011001100110011001100110",
18826 => "011001100110011001100110",
18827 => "011101100110001000100011",
18828 => "011111110110000000000000",
18829 => "010101110100001000000000",
18830 => "000000000000000000000000",
18831 => "000000000000000000000000",
18832 => "010000110100001101000011",
18833 => "010000110100001101000011",
18834 => "010000110100001101000011",
18835 => "010000110100001101000011",
18836 => "010000110100001101000011",
18837 => "010000110100001101000011",
18838 => "010000110100001101000011",
18839 => "010000110100001101000011",
18840 => "010000110100001101000011",
18841 => "010000110100001101000011",
18842 => "010000110100001101000011",
18843 => "001100100011001000110010",
18844 => "000000000000000000000000",
18845 => "000000000000000000000000",
18846 => "000000000000000000000000",
18847 => "000000000000000000000000",
18848 => "000000000000000000000000",
18849 => "000000000000000000000000",
18850 => "000000000000000000000000",
18851 => "000000000000000000000000",
18852 => "000000000000000000000000",
18853 => "000000000000000000000000",
18854 => "000000000000000000000000",
18855 => "000000000000000000000000",
18856 => "000000000000000000000000",
18857 => "000000000000000000000000",
18858 => "000000000000000000000000",
18859 => "000000000000000000000000",
18860 => "000000000000000000000000",
18861 => "000000000000000000000000",
18862 => "000000000000000000000000",
18863 => "000000000000000000000000",
18864 => "000000000000000000000000",
18865 => "000000000000000000000000",
18866 => "000000000000000000000000",
18867 => "000000000000000000000000",
18868 => "000000000000000000000000",
18869 => "000000000000000000000000",
18870 => "000000000000000000000000",
18871 => "000000000000000000000000",
18872 => "000000000000000000000000",
18873 => "000000000000000000000000",
18874 => "000000000000000000000000",
18875 => "000000000000000000000000",
18876 => "000000000000000000000000",
18877 => "000000000000000000000000",
18878 => "000000000000000000000000",
18879 => "000000000000000000000000",
18880 => "000000000000000000000000",
18881 => "000000000000000000000000",
18882 => "000000000000000000000000",
18883 => "000000000000000000000000",
18884 => "000000000000000000000000",
18885 => "000000000000000000000000",
18886 => "000000000000000000000000",
18887 => "000000000000000000000000",
18888 => "000000000000000000000000",
18889 => "000000000000000000000000",
18890 => "000000000000000000000000",
18891 => "000000000000000000000000",
18892 => "000000000000000000000000",
18893 => "000000000000000000000000",
18894 => "000000000000000000000000",
18895 => "000000000000000000000000",
18896 => "000000000000000000000000",
18897 => "000000000000000000000000",
18898 => "000000000000000000000000",
18899 => "000000000000000000000000",
18900 => "000000000000000000000000",
18901 => "000000000000000000000000",
18902 => "000000000000000000000000",
18903 => "000000000000000000000000",
18904 => "000000000000000000000000",
18905 => "000000000000000000000000",
18906 => "000000000000000000000000",
18907 => "000000000000000000000000",
18908 => "000000000000000000000000",
18909 => "000000000000000000000000",
18910 => "000000000000000000000000",
18911 => "000000000000000000000000",
18912 => "000000000000000000000000",
18913 => "000000000000000000000000",
18914 => "000000000000000000000000",
18915 => "000000000000000000000000",
18916 => "000000000000000000000000",
18917 => "000000000000000000000000",
18918 => "000000000000000000000000",
18919 => "000000000000000000000000",
18920 => "000000000000000000000000",
18921 => "000000000000000000000000",
18922 => "000000000000000000000000",
18923 => "000000000000000000000000",
18924 => "000000000000000000000000",
18925 => "000000000000000000000000",
18926 => "000000000000000000000000",
18927 => "000000000000000000000000",
18928 => "000000000000000000000000",
18929 => "000000000000000000000000",
18930 => "000000000000000000000000",
18931 => "000000000000000000000000",
18932 => "000000000000000000000000",
18933 => "000000000000000000000000",
18934 => "000000000000000000000000",
18935 => "000000000000000000000000",
18936 => "000000000000000000000000",
18937 => "000000000000000000000000",
18938 => "000000000000000000000000",
18939 => "000000000000000000000000",
18940 => "000000000000000000000000",
18941 => "000000000000000000000000",
18942 => "000110100001101000011010",
18943 => "000111010001110100011101",
18944 => "001011110010111100101111",
18945 => "010000110100001101000011",
18946 => "010000110100001101000011",
18947 => "010000110100001101000011",
18948 => "010000110100001101000011",
18949 => "010000110100001101000011",
18950 => "010000110100001101000011",
18951 => "010000110100001101000011",
18952 => "010000110100001101000011",
18953 => "010000110100001101000011",
18954 => "010000110100001101000011",
18955 => "010000110100001101000011",
18956 => "000011100000111000001110",
18957 => "000000000000000000000000",
18958 => "001101000010011100000000",
18959 => "011111110110000000000000",
18960 => "011111010110000000000110",
18961 => "011001100110011001100110",
18962 => "011001100110011001100110",
18963 => "011110000110001000011100",
18964 => "011111110110000000000000",
18965 => "011101100110001000100110",
18966 => "011001100110011001100110",
18967 => "011000110110001101100011",
18968 => "000000000000000000000000",
18969 => "000000000000000000000000",
18970 => "010001100100011001000110",
18971 => "011001100110011001100110",
18972 => "011011110110010001000011",
18973 => "011111110110000000000000",
18974 => "011111110110000000000000",
18975 => "011001100110011001100110",
18976 => "011001100110011001100110",
18977 => "011101100110001000100011",
18978 => "011111110110000000000000",
18979 => "010101110100001000000000",
18980 => "000000000000000000000000",
18981 => "000000000000000000000000",
18982 => "010000110100001101000011",
18983 => "010000110100001101000011",
18984 => "010000110100001101000011",
18985 => "010000110100001101000011",
18986 => "010000110100001101000011",
18987 => "010000110100001101000011",
18988 => "010000110100001101000011",
18989 => "010000110100001101000011",
18990 => "010000110100001101000011",
18991 => "010000110100001101000011",
18992 => "010000110100001101000011",
18993 => "001110100011101000111010",
18994 => "000111010001110100011101",
18995 => "000111010001110100011101",
18996 => "000000010000000100000001",
18997 => "000000000000000000000000",
18998 => "000000000000000000000000",
18999 => "000000000000000000000000",
19000 => "000000000000000000000000",
19001 => "000000000000000000000000",
19002 => "000000000000000000000000",
19003 => "000000000000000000000000",
19004 => "000000000000000000000000",
19005 => "000000000000000000000000",
19006 => "000000000000000000000000",
19007 => "000000000000000000000000",
19008 => "000000000000000000000000",
19009 => "000000000000000000000000",
19010 => "000000000000000000000000",
19011 => "000000000000000000000000",
19012 => "000000000000000000000000",
19013 => "000000000000000000000000",
19014 => "000000000000000000000000",
19015 => "000000000000000000000000",
19016 => "000000000000000000000000",
19017 => "000000000000000000000000",
19018 => "000000000000000000000000",
19019 => "000000000000000000000000",
19020 => "000000000000000000000000",
19021 => "000000000000000000000000",
19022 => "000000000000000000000000",
19023 => "000000000000000000000000",
19024 => "000000000000000000000000",
19025 => "000000000000000000000000",
19026 => "000000000000000000000000",
19027 => "000000000000000000000000",
19028 => "000000000000000000000000",
19029 => "000000000000000000000000",
19030 => "000000000000000000000000",
19031 => "000000000000000000000000",
19032 => "000000000000000000000000",
19033 => "000000000000000000000000",
19034 => "000000000000000000000000",
19035 => "000000000000000000000000",
19036 => "000000000000000000000000",
19037 => "000000000000000000000000",
19038 => "000000000000000000000000",
19039 => "000000000000000000000000",
19040 => "000000000000000000000000",
19041 => "000000000000000000000000",
19042 => "000000000000000000000000",
19043 => "000000000000000000000000",
19044 => "000000000000000000000000",
19045 => "000000000000000000000000",
19046 => "000000000000000000000000",
19047 => "000000000000000000000000",
19048 => "000000000000000000000000",
19049 => "000000000000000000000000",
19050 => "000000000000000000000000",
19051 => "000000000000000000000000",
19052 => "000000000000000000000000",
19053 => "000000000000000000000000",
19054 => "000000000000000000000000",
19055 => "000000000000000000000000",
19056 => "000000000000000000000000",
19057 => "000000000000000000000000",
19058 => "000000000000000000000000",
19059 => "000000000000000000000000",
19060 => "000000000000000000000000",
19061 => "000000000000000000000000",
19062 => "000000000000000000000000",
19063 => "000000000000000000000000",
19064 => "000000000000000000000000",
19065 => "000000000000000000000000",
19066 => "000000000000000000000000",
19067 => "000000000000000000000000",
19068 => "000000000000000000000000",
19069 => "000000000000000000000000",
19070 => "000000000000000000000000",
19071 => "000000000000000000000000",
19072 => "000000000000000000000000",
19073 => "000000000000000000000000",
19074 => "000000000000000000000000",
19075 => "000000000000000000000000",
19076 => "000000000000000000000000",
19077 => "000000000000000000000000",
19078 => "000000000000000000000000",
19079 => "000000000000000000000000",
19080 => "000000000000000000000000",
19081 => "000000000000000000000000",
19082 => "000000000000000000000000",
19083 => "000000000000000000000000",
19084 => "000000000000000000000000",
19085 => "000000000000000000000000",
19086 => "000000000000000000000000",
19087 => "000000000000000000000000",
19088 => "000000000000000000000000",
19089 => "000000000000000000000000",
19090 => "000000000000000000000000",
19091 => "000000000000000000000000",
19092 => "001110110011101100111011",
19093 => "010000110100001101000011",
19094 => "010000110100001101000011",
19095 => "010000110100001101000011",
19096 => "010000110100001101000011",
19097 => "010000110100001101000011",
19098 => "010000110100001101000011",
19099 => "010000110100001101000011",
19100 => "010000110100001101000011",
19101 => "010000110100001101000011",
19102 => "010000110100001101000011",
19103 => "010000110100001101000011",
19104 => "010000110100001101000011",
19105 => "010000110100001101000011",
19106 => "000011100000111000001110",
19107 => "000000000000000000000000",
19108 => "001101000010011100000000",
19109 => "011111110110000000000000",
19110 => "011111010110000000000110",
19111 => "011001100110011001100110",
19112 => "011001100110011001100110",
19113 => "011110000110001000011100",
19114 => "011111110110000000000000",
19115 => "011101100110001000100110",
19116 => "011001100110011001100110",
19117 => "011000110110001101100011",
19118 => "000000000000000000000000",
19119 => "000000000000000000000000",
19120 => "010001100100011001000110",
19121 => "011001100110011001100110",
19122 => "011011110110010001000011",
19123 => "011111110110000000000000",
19124 => "011111110110000000000000",
19125 => "011001100110011001100110",
19126 => "011001100110011001100110",
19127 => "011101100110001000100011",
19128 => "011111110110000000000000",
19129 => "010101110100001000000000",
19130 => "000000000000000000000000",
19131 => "000000000000000000000000",
19132 => "010000110100001101000011",
19133 => "010000110100001101000011",
19134 => "010000110100001101000011",
19135 => "010000110100001101000011",
19136 => "010000110100001101000011",
19137 => "010000110100001101000011",
19138 => "010000110100001101000011",
19139 => "010000110100001101000011",
19140 => "010000110100001101000011",
19141 => "010000110100001101000011",
19142 => "010000110100001101000011",
19143 => "010000110100001101000011",
19144 => "010000110100001101000011",
19145 => "010000110100001101000011",
19146 => "000000100000001000000010",
19147 => "000000000000000000000000",
19148 => "000000000000000000000000",
19149 => "000000000000000000000000",
19150 => "000000000000000000000000",
19151 => "000000000000000000000000",
19152 => "000000000000000000000000",
19153 => "000000000000000000000000",
19154 => "000000000000000000000000",
19155 => "000000000000000000000000",
19156 => "000000000000000000000000",
19157 => "000000000000000000000000",
19158 => "000000000000000000000000",
19159 => "000000000000000000000000",
19160 => "000000000000000000000000",
19161 => "000000000000000000000000",
19162 => "000000000000000000000000",
19163 => "000000000000000000000000",
19164 => "000000000000000000000000",
19165 => "000000000000000000000000",
19166 => "000000000000000000000000",
19167 => "000000000000000000000000",
19168 => "000000000000000000000000",
19169 => "000000000000000000000000",
19170 => "000000000000000000000000",
19171 => "000000000000000000000000",
19172 => "000000000000000000000000",
19173 => "000000000000000000000000",
19174 => "000000000000000000000000",
19175 => "000000000000000000000000",
19176 => "000000000000000000000000",
19177 => "000000000000000000000000",
19178 => "000000000000000000000000",
19179 => "000000000000000000000000",
19180 => "000000000000000000000000",
19181 => "000000000000000000000000",
19182 => "000000000000000000000000",
19183 => "000000000000000000000000",
19184 => "000000000000000000000000",
19185 => "000000000000000000000000",
19186 => "000000000000000000000000",
19187 => "000000000000000000000000",
19188 => "000000000000000000000000",
19189 => "000000000000000000000000",
19190 => "000000000000000000000000",
19191 => "000000000000000000000000",
19192 => "000000000000000000000000",
19193 => "000000000000000000000000",
19194 => "000000000000000000000000",
19195 => "000000000000000000000000",
19196 => "000000000000000000000000",
19197 => "000000000000000000000000",
19198 => "000000000000000000000000",
19199 => "000000000000000000000000",
19200 => "000000000000000000000000",
19201 => "000000000000000000000000",
19202 => "000000000000000000000000",
19203 => "000000000000000000000000",
19204 => "000000000000000000000000",
19205 => "000000000000000000000000",
19206 => "000000000000000000000000",
19207 => "000000000000000000000000",
19208 => "000000000000000000000000",
19209 => "000000000000000000000000",
19210 => "000000000000000000000000",
19211 => "000000000000000000000000",
19212 => "000000000000000000000000",
19213 => "000000000000000000000000",
19214 => "000000000000000000000000",
19215 => "000000000000000000000000",
19216 => "000000000000000000000000",
19217 => "000000000000000000000000",
19218 => "000000000000000000000000",
19219 => "000000000000000000000000",
19220 => "000000000000000000000000",
19221 => "000000000000000000000000",
19222 => "000000000000000000000000",
19223 => "000000000000000000000000",
19224 => "000000000000000000000000",
19225 => "000000000000000000000000",
19226 => "000000000000000000000000",
19227 => "000000000000000000000000",
19228 => "000000000000000000000000",
19229 => "000000000000000000000000",
19230 => "000000000000000000000000",
19231 => "000000000000000000000000",
19232 => "000000000000000000000000",
19233 => "000000000000000000000000",
19234 => "000000000000000000000000",
19235 => "000000000000000000000000",
19236 => "000000000000000000000000",
19237 => "000000000000000000000000",
19238 => "000000000000000000000000",
19239 => "000000010000000100000001",
19240 => "000010100000101000001010",
19241 => "000010100000101000001010",
19242 => "001111000011110000111100",
19243 => "010000110100001101000011",
19244 => "010000110100001101000011",
19245 => "010000110100001101000011",
19246 => "010000110100001101000011",
19247 => "010000110100001101000011",
19248 => "010000110100001101000011",
19249 => "010000110100001101000011",
19250 => "010000110100001101000011",
19251 => "010000110100001101000011",
19252 => "010000110100001101000011",
19253 => "010000110100001101000011",
19254 => "010000110100001101000011",
19255 => "010000110100001101000011",
19256 => "000011100000111000001110",
19257 => "000000000000000000000000",
19258 => "001101000010011100000000",
19259 => "011111110110000000000000",
19260 => "011111010110000000000110",
19261 => "011001100110011001100110",
19262 => "011001100110011001100110",
19263 => "011110000110001000011100",
19264 => "011111110110000000000000",
19265 => "011101100110001000100110",
19266 => "011001100110011001100110",
19267 => "011000110110001101100011",
19268 => "000000000000000000000000",
19269 => "000000000000000000000000",
19270 => "010001100100011001000110",
19271 => "011001100110011001100110",
19272 => "011011110110010001000011",
19273 => "011111110110000000000000",
19274 => "011111110110000000000000",
19275 => "011001100110011001100110",
19276 => "011001100110011001100110",
19277 => "011101100110001000100011",
19278 => "011111110110000000000000",
19279 => "010101110100001000000000",
19280 => "000000000000000000000000",
19281 => "000000000000000000000000",
19282 => "010000110100001101000011",
19283 => "010000110100001101000011",
19284 => "010000110100001101000011",
19285 => "010000110100001101000011",
19286 => "010000110100001101000011",
19287 => "010000110100001101000011",
19288 => "010000110100001101000011",
19289 => "010000110100001101000011",
19290 => "010000110100001101000011",
19291 => "010000110100001101000011",
19292 => "010000110100001101000011",
19293 => "010001000100010001000100",
19294 => "010001100100011001000110",
19295 => "010001100100011001000110",
19296 => "000010000000100000001000",
19297 => "000001100000011000000110",
19298 => "000000110000001100000011",
19299 => "000000000000000000000000",
19300 => "000000000000000000000000",
19301 => "000000000000000000000000",
19302 => "000000000000000000000000",
19303 => "000000000000000000000000",
19304 => "000000000000000000000000",
19305 => "000000000000000000000000",
19306 => "000000000000000000000000",
19307 => "000000000000000000000000",
19308 => "000000000000000000000000",
19309 => "000000000000000000000000",
19310 => "000000000000000000000000",
19311 => "000000000000000000000000",
19312 => "000000000000000000000000",
19313 => "000000000000000000000000",
19314 => "000000000000000000000000",
19315 => "000000000000000000000000",
19316 => "000000000000000000000000",
19317 => "000000000000000000000000",
19318 => "000000000000000000000000",
19319 => "000000000000000000000000",
19320 => "000000000000000000000000",
19321 => "000000000000000000000000",
19322 => "000000000000000000000000",
19323 => "000000000000000000000000",
19324 => "000000000000000000000000",
19325 => "000000000000000000000000",
19326 => "000000000000000000000000",
19327 => "000000000000000000000000",
19328 => "000000000000000000000000",
19329 => "000000000000000000000000",
19330 => "000000000000000000000000",
19331 => "000000000000000000000000",
19332 => "000000000000000000000000",
19333 => "000000000000000000000000",
19334 => "000000000000000000000000",
19335 => "000000000000000000000000",
19336 => "000000000000000000000000",
19337 => "000000000000000000000000",
19338 => "000000000000000000000000",
19339 => "000000000000000000000000",
19340 => "000000000000000000000000",
19341 => "000000000000000000000000",
19342 => "000000000000000000000000",
19343 => "000000000000000000000000",
19344 => "000000000000000000000000",
19345 => "000000000000000000000000",
19346 => "000000000000000000000000",
19347 => "000000000000000000000000",
19348 => "000000000000000000000000",
19349 => "000000000000000000000000",
19350 => "000000000000000000000000",
19351 => "000000000000000000000000",
19352 => "000000000000000000000000",
19353 => "000000000000000000000000",
19354 => "000000000000000000000000",
19355 => "000000000000000000000000",
19356 => "000000000000000000000000",
19357 => "000000000000000000000000",
19358 => "000000000000000000000000",
19359 => "000000000000000000000000",
19360 => "000000000000000000000000",
19361 => "000000000000000000000000",
19362 => "000000000000000000000000",
19363 => "000000000000000000000000",
19364 => "000000000000000000000000",
19365 => "000000000000000000000000",
19366 => "000000000000000000000000",
19367 => "000000000000000000000000",
19368 => "000000000000000000000000",
19369 => "000000000000000000000000",
19370 => "000000000000000000000000",
19371 => "000000000000000000000000",
19372 => "000000000000000000000000",
19373 => "000000000000000000000000",
19374 => "000000000000000000000000",
19375 => "000000000000000000000000",
19376 => "000000000000000000000000",
19377 => "000000000000000000000000",
19378 => "000000000000000000000000",
19379 => "000000000000000000000000",
19380 => "000000000000000000000000",
19381 => "000000000000000000000000",
19382 => "000000000000000000000000",
19383 => "000000000000000000000000",
19384 => "000000000000000000000000",
19385 => "000000000000000000000000",
19386 => "000000000000000000000000",
19387 => "000000000000000000000000",
19388 => "000000000000000000000000",
19389 => "000100000001000000010000",
19390 => "011001100110011001100110",
19391 => "011001100110011001100110",
19392 => "010001110100011101000111",
19393 => "010000110100001101000011",
19394 => "010000110100001101000011",
19395 => "010000110100001101000011",
19396 => "010000110100001101000011",
19397 => "010000110100001101000011",
19398 => "010000110100001101000011",
19399 => "010000110100001101000011",
19400 => "010000110100001101000011",
19401 => "010000110100001101000011",
19402 => "010000110100001101000011",
19403 => "010000110100001101000011",
19404 => "010000110100001101000011",
19405 => "010000110100001101000011",
19406 => "000011100000111000001110",
19407 => "000000000000000000000000",
19408 => "001101000010011100000000",
19409 => "011111110110000000000000",
19410 => "011111010110000000000110",
19411 => "011001100110011001100110",
19412 => "011001100110011001100110",
19413 => "011110000110001000011100",
19414 => "011111110110000000000000",
19415 => "011101100110001000100110",
19416 => "011001100110011001100110",
19417 => "011000110110001101100011",
19418 => "000000000000000000000000",
19419 => "000000000000000000000000",
19420 => "010001100100011001000110",
19421 => "011001100110011001100110",
19422 => "011011110110010001000011",
19423 => "011111110110000000000000",
19424 => "011111110110000000000000",
19425 => "011001100110011001100110",
19426 => "011001100110011001100110",
19427 => "011101100110001000100011",
19428 => "011111110110000000000000",
19429 => "010101110100001000000000",
19430 => "000000000000000000000000",
19431 => "000000000000000000000000",
19432 => "010000110100001101000011",
19433 => "010000110100001101000011",
19434 => "010000110100001101000011",
19435 => "010000110100001101000011",
19436 => "010000110100001101000011",
19437 => "010000110100001101000011",
19438 => "010000110100001101000011",
19439 => "010000110100001101000011",
19440 => "010000110100001101000011",
19441 => "010000110100001101000011",
19442 => "010000110100001101000011",
19443 => "010011000100110001001100",
19444 => "011001100110011001100110",
19445 => "011001100110011001100110",
19446 => "010001000100010001000100",
19447 => "010000110100001101000011",
19448 => "000111010001110100011101",
19449 => "000000000000000000000000",
19450 => "000000000000000000000000",
19451 => "000000000000000000000000",
19452 => "000000000000000000000000",
19453 => "000000000000000000000000",
19454 => "000000000000000000000000",
19455 => "000000000000000000000000",
19456 => "000000000000000000000000",
19457 => "000000000000000000000000",
19458 => "000000000000000000000000",
19459 => "000000000000000000000000",
19460 => "000000000000000000000000",
19461 => "000000000000000000000000",
19462 => "000000000000000000000000",
19463 => "000000000000000000000000",
19464 => "000000000000000000000000",
19465 => "000000000000000000000000",
19466 => "000000000000000000000000",
19467 => "000000000000000000000000",
19468 => "000000000000000000000000",
19469 => "000000000000000000000000",
19470 => "000000000000000000000000",
19471 => "000000000000000000000000",
19472 => "000000000000000000000000",
19473 => "000000000000000000000000",
19474 => "000000000000000000000000",
19475 => "000000000000000000000000",
19476 => "000000000000000000000000",
19477 => "000000000000000000000000",
19478 => "000000000000000000000000",
19479 => "000000000000000000000000",
19480 => "000000000000000000000000",
19481 => "000000000000000000000000",
19482 => "000000000000000000000000",
19483 => "000000000000000000000000",
19484 => "000000000000000000000000",
19485 => "000000000000000000000000",
19486 => "000000000000000000000000",
19487 => "000000000000000000000000",
19488 => "000000000000000000000000",
19489 => "000000000000000000000000",
19490 => "000000000000000000000000",
19491 => "000000000000000000000000",
19492 => "000000000000000000000000",
19493 => "000000000000000000000000",
19494 => "000000000000000000000000",
19495 => "000000000000000000000000",
19496 => "000000000000000000000000",
19497 => "000000000000000000000000",
19498 => "000000000000000000000000",
19499 => "000000000000000000000000",
19500 => "000000000000000000000000",
19501 => "000000000000000000000000",
19502 => "000000000000000000000000",
19503 => "000000000000000000000000",
19504 => "000000000000000000000000",
19505 => "000000000000000000000000",
19506 => "000000000000000000000000",
19507 => "000000000000000000000000",
19508 => "000000000000000000000000",
19509 => "000000000000000000000000",
19510 => "000000000000000000000000",
19511 => "000000000000000000000000",
19512 => "000000000000000000000000",
19513 => "000000000000000000000000",
19514 => "000000000000000000000000",
19515 => "000000000000000000000000",
19516 => "000000000000000000000000",
19517 => "000000000000000000000000",
19518 => "000000000000000000000000",
19519 => "000000000000000000000000",
19520 => "000000000000000000000000",
19521 => "000000000000000000000000",
19522 => "000000000000000000000000",
19523 => "000000000000000000000000",
19524 => "000000000000000000000000",
19525 => "000000000000000000000000",
19526 => "000000000000000000000000",
19527 => "000000000000000000000000",
19528 => "000000000000000000000000",
19529 => "000000000000000000000000",
19530 => "000000000000000000000000",
19531 => "000000000000000000000000",
19532 => "000000000000000000000000",
19533 => "000000000000000000000000",
19534 => "000000000000000000000000",
19535 => "000000000000000000000000",
19536 => "000000000000000000000000",
19537 => "000000000000000000000000",
19538 => "000000000000000000000000",
19539 => "000100000001000000010000",
19540 => "011001100110011001100110",
19541 => "011001100110011001100110",
19542 => "010001110100011101000111",
19543 => "010000110100001101000011",
19544 => "010000110100001101000011",
19545 => "010000110100001101000011",
19546 => "010000110100001101000011",
19547 => "010000110100001101000011",
19548 => "010000110100001101000011",
19549 => "010000110100001101000011",
19550 => "010000110100001101000011",
19551 => "010000110100001101000011",
19552 => "010000110100001101000011",
19553 => "010000110100001101000011",
19554 => "010000110100001101000011",
19555 => "010000110100001101000011",
19556 => "000011100000111000001110",
19557 => "000000000000000000000000",
19558 => "001101000010011100000000",
19559 => "011111110110000000000000",
19560 => "011111010110000000000110",
19561 => "011001100110011001100110",
19562 => "011001100110011001100110",
19563 => "011110000110001000011100",
19564 => "011111110110000000000000",
19565 => "011101100110001000100110",
19566 => "011001100110011001100110",
19567 => "011000110110001101100011",
19568 => "000000000000000000000000",
19569 => "000000000000000000000000",
19570 => "010001100100011001000110",
19571 => "011001100110011001100110",
19572 => "011011110110010001000011",
19573 => "011111110110000000000000",
19574 => "011111110110000000000000",
19575 => "011001100110011001100110",
19576 => "011001100110011001100110",
19577 => "011101100110001000100011",
19578 => "011111110110000000000000",
19579 => "010101110100001000000000",
19580 => "000000000000000000000000",
19581 => "000000000000000000000000",
19582 => "010000110100001101000011",
19583 => "010000110100001101000011",
19584 => "010000110100001101000011",
19585 => "010000110100001101000011",
19586 => "010000110100001101000011",
19587 => "010000110100001101000011",
19588 => "010000110100001101000011",
19589 => "010000110100001101000011",
19590 => "010000110100001101000011",
19591 => "010000110100001101000011",
19592 => "010000110100001101000011",
19593 => "010011000100110001001100",
19594 => "011001100110011001100110",
19595 => "011001100110011001100110",
19596 => "010001000100010001000100",
19597 => "010000110100001101000011",
19598 => "000111010001110100011101",
19599 => "000000000000000000000000",
19600 => "000000000000000000000000",
19601 => "000000000000000000000000",
19602 => "000000000000000000000000",
19603 => "000000000000000000000000",
19604 => "000000000000000000000000",
19605 => "000000000000000000000000",
19606 => "000000000000000000000000",
19607 => "000000000000000000000000",
19608 => "000000000000000000000000",
19609 => "000000000000000000000000",
19610 => "000000000000000000000000",
19611 => "000000000000000000000000",
19612 => "000000000000000000000000",
19613 => "000000000000000000000000",
19614 => "000000000000000000000000",
19615 => "000000000000000000000000",
19616 => "000000000000000000000000",
19617 => "000000000000000000000000",
19618 => "000000000000000000000000",
19619 => "000000000000000000000000",
19620 => "000000000000000000000000",
19621 => "000000000000000000000000",
19622 => "000000000000000000000000",
19623 => "000000000000000000000000",
19624 => "000000000000000000000000",
19625 => "000000000000000000000000",
19626 => "000000000000000000000000",
19627 => "000000000000000000000000",
19628 => "000000000000000000000000",
19629 => "000000000000000000000000",
19630 => "000000000000000000000000",
19631 => "000000000000000000000000",
19632 => "000000000000000000000000",
19633 => "000000000000000000000000",
19634 => "000000000000000000000000",
19635 => "000000000000000000000000",
19636 => "000000000000000000000000",
19637 => "000000000000000000000000",
19638 => "000000000000000000000000",
19639 => "000000000000000000000000",
19640 => "000000000000000000000000",
19641 => "000000000000000000000000",
19642 => "000000000000000000000000",
19643 => "000000000000000000000000",
19644 => "000000000000000000000000",
19645 => "000000000000000000000000",
19646 => "000000000000000000000000",
19647 => "000000000000000000000000",
19648 => "000000000000000000000000",
19649 => "000000000000000000000000",
19650 => "000000000000000000000000",
19651 => "000000000000000000000000",
19652 => "000000000000000000000000",
19653 => "000000000000000000000000",
19654 => "000000000000000000000000",
19655 => "000000000000000000000000",
19656 => "000000000000000000000000",
19657 => "000000000000000000000000",
19658 => "000000000000000000000000",
19659 => "000000000000000000000000",
19660 => "000000000000000000000000",
19661 => "000000000000000000000000",
19662 => "000000000000000000000000",
19663 => "000000000000000000000000",
19664 => "000000000000000000000000",
19665 => "000000000000000000000000",
19666 => "000000000000000000000000",
19667 => "000000000000000000000000",
19668 => "000000000000000000000000",
19669 => "000000000000000000000000",
19670 => "000000000000000000000000",
19671 => "000000000000000000000000",
19672 => "000000000000000000000000",
19673 => "000000000000000000000000",
19674 => "000000000000000000000000",
19675 => "000000000000000000000000",
19676 => "000000000000000000000000",
19677 => "000000000000000000000000",
19678 => "000000000000000000000000",
19679 => "000000000000000000000000",
19680 => "000000000000000000000000",
19681 => "000000000000000000000000",
19682 => "000000000000000000000000",
19683 => "000000000000000000000000",
19684 => "000000000000000000000000",
19685 => "000000000000000000000000",
19686 => "000000000000000000000000",
19687 => "000110100001101000011010",
19688 => "001101010011010100110101",
19689 => "001111000011110000111100",
19690 => "011001100110011001100110",
19691 => "011001100110011001100110",
19692 => "010001110100011101000111",
19693 => "010000110100001101000011",
19694 => "010000110100001101000011",
19695 => "010000110100001101000011",
19696 => "010000110100001101000011",
19697 => "010000110100001101000011",
19698 => "010000110100001101000011",
19699 => "010000110100001101000011",
19700 => "010000110100001101000011",
19701 => "010000110100001101000011",
19702 => "010000110100001101000011",
19703 => "001111100011111000111110",
19704 => "000011100000111000001110",
19705 => "000011100000111000001110",
19706 => "000000110000001100000011",
19707 => "000000000000000000000000",
19708 => "000010110000100000000000",
19709 => "000110110001010000000000",
19710 => "001000000001101000000110",
19711 => "011001100110011001100110",
19712 => "011001100110011001100110",
19713 => "011010100110010101010110",
19714 => "011010110110010101010000",
19715 => "010010110100011100111010",
19716 => "000101100001011000010110",
19717 => "000101010001010100010101",
19718 => "000000000000000000000000",
19719 => "000000000000000000000000",
19720 => "000011110000111100001111",
19721 => "000101100001011000010110",
19722 => "001100110011000100101010",
19723 => "011010110110010101010000",
19724 => "011010110110010101010000",
19725 => "011001100110011001100110",
19726 => "011001100110011001100110",
19727 => "001101010011000100100011",
19728 => "000110110001010000000000",
19729 => "000100110000111000000000",
19730 => "000000000000000000000000",
19731 => "000000000000000000000000",
19732 => "000011100000111000001110",
19733 => "000011100000111000001110",
19734 => "001011110010111100101111",
19735 => "010000110100001101000011",
19736 => "010000110100001101000011",
19737 => "010000110100001101000011",
19738 => "010000110100001101000011",
19739 => "010000110100001101000011",
19740 => "010000110100001101000011",
19741 => "010000110100001101000011",
19742 => "010000110100001101000011",
19743 => "010011000100110001001100",
19744 => "011001100110011001100110",
19745 => "011001100110011001100110",
19746 => "010001000100010001000100",
19747 => "010000110100001101000011",
19748 => "001110110011101100111011",
19749 => "001101010011010100110101",
19750 => "001010010010100100101001",
19751 => "000000000000000000000000",
19752 => "000000000000000000000000",
19753 => "000000000000000000000000",
19754 => "000000000000000000000000",
19755 => "000000000000000000000000",
19756 => "000000000000000000000000",
19757 => "000000000000000000000000",
19758 => "000000000000000000000000",
19759 => "000000000000000000000000",
19760 => "000000000000000000000000",
19761 => "000000000000000000000000",
19762 => "000000000000000000000000",
19763 => "000000000000000000000000",
19764 => "000000000000000000000000",
19765 => "000000000000000000000000",
19766 => "000000000000000000000000",
19767 => "000000000000000000000000",
19768 => "000000000000000000000000",
19769 => "000000000000000000000000",
19770 => "000000000000000000000000",
19771 => "000000000000000000000000",
19772 => "000000000000000000000000",
19773 => "000000000000000000000000",
19774 => "000000000000000000000000",
19775 => "000000000000000000000000",
19776 => "000000000000000000000000",
19777 => "000000000000000000000000",
19778 => "000000000000000000000000",
19779 => "000000000000000000000000",
19780 => "000000000000000000000000",
19781 => "000000000000000000000000",
19782 => "000000000000000000000000",
19783 => "000000000000000000000000",
19784 => "000000000000000000000000",
19785 => "000000000000000000000000",
19786 => "000000000000000000000000",
19787 => "000000000000000000000000",
19788 => "000000000000000000000000",
19789 => "000000000000000000000000",
19790 => "000000000000000000000000",
19791 => "000000000000000000000000",
19792 => "000000000000000000000000",
19793 => "000000000000000000000000",
19794 => "000000000000000000000000",
19795 => "000000000000000000000000",
19796 => "000000000000000000000000",
19797 => "000000000000000000000000",
19798 => "000000000000000000000000",
19799 => "000000000000000000000000",
19800 => "000000000000000000000000",
19801 => "000000000000000000000000",
19802 => "000000000000000000000000",
19803 => "000000000000000000000000",
19804 => "000000000000000000000000",
19805 => "000000000000000000000000",
19806 => "000000000000000000000000",
19807 => "000000000000000000000000",
19808 => "000000000000000000000000",
19809 => "000000000000000000000000",
19810 => "000000000000000000000000",
19811 => "000000000000000000000000",
19812 => "000000000000000000000000",
19813 => "000000000000000000000000",
19814 => "000000000000000000000000",
19815 => "000000000000000000000000",
19816 => "000000000000000000000000",
19817 => "000000000000000000000000",
19818 => "000000000000000000000000",
19819 => "000000000000000000000000",
19820 => "000000000000000000000000",
19821 => "000000000000000000000000",
19822 => "000000000000000000000000",
19823 => "000000000000000000000000",
19824 => "000000000000000000000000",
19825 => "000000000000000000000000",
19826 => "000000000000000000000000",
19827 => "000000000000000000000000",
19828 => "000000000000000000000000",
19829 => "000000000000000000000000",
19830 => "000000000000000000000000",
19831 => "000000000000000000000000",
19832 => "000000000000000000000000",
19833 => "000000000000000000000000",
19834 => "000000000000000000000000",
19835 => "000000000000000000000000",
19836 => "000000000000000000000000",
19837 => "001000100010001000100010",
19838 => "010000110100001101000011",
19839 => "010010000100100001001000",
19840 => "011001100110011001100110",
19841 => "011001100110011001100110",
19842 => "010001110100011101000111",
19843 => "010000110100001101000011",
19844 => "010000110100001101000011",
19845 => "010000110100001101000011",
19846 => "010000110100001101000011",
19847 => "010000110100001101000011",
19848 => "010000110100001101000011",
19849 => "010000110100001101000011",
19850 => "010000110100001101000011",
19851 => "010000110100001101000011",
19852 => "010000110100001101000011",
19853 => "001111010011110100111101",
19854 => "000000000000000000000000",
19855 => "000000000000000000000000",
19856 => "000000000000000000000000",
19857 => "000000000000000000000000",
19858 => "000000000000000000000000",
19859 => "000000000000000000000000",
19860 => "000001100000011000000110",
19861 => "011001100110011001100110",
19862 => "011001100110011001100110",
19863 => "011001100110011001100110",
19864 => "011001100110011001100110",
19865 => "010000000100000001000000",
19866 => "000000000000000000000000",
19867 => "000000000000000000000000",
19868 => "000000000000000000000000",
19869 => "000000000000000000000000",
19870 => "000000000000000000000000",
19871 => "000000000000000000000000",
19872 => "001000110010001100100011",
19873 => "011001100110011001100110",
19874 => "011001100110011001100110",
19875 => "011001100110011001100110",
19876 => "011001100110011001100110",
19877 => "001000110010001100100011",
19878 => "000000000000000000000000",
19879 => "000000000000000000000000",
19880 => "000000000000000000000000",
19881 => "000000000000000000000000",
19882 => "000000000000000000000000",
19883 => "000000000000000000000000",
19884 => "001010100010101000101010",
19885 => "010000110100001101000011",
19886 => "010000110100001101000011",
19887 => "010000110100001101000011",
19888 => "010000110100001101000011",
19889 => "010000110100001101000011",
19890 => "010000110100001101000011",
19891 => "010000110100001101000011",
19892 => "010000110100001101000011",
19893 => "010011000100110001001100",
19894 => "011001100110011001100110",
19895 => "011001100110011001100110",
19896 => "010001000100010001000100",
19897 => "010000110100001101000011",
19898 => "010000110100001101000011",
19899 => "010000110100001101000011",
19900 => "001101000011010000110100",
19901 => "000000000000000000000000",
19902 => "000000000000000000000000",
19903 => "000000000000000000000000",
19904 => "000000000000000000000000",
19905 => "000000000000000000000000",
19906 => "000000000000000000000000",
19907 => "000000000000000000000000",
19908 => "000000000000000000000000",
19909 => "000000000000000000000000",
19910 => "000000000000000000000000",
19911 => "000000000000000000000000",
19912 => "000000000000000000000000",
19913 => "000000000000000000000000",
19914 => "000000000000000000000000",
19915 => "000000000000000000000000",
19916 => "000000000000000000000000",
19917 => "000000000000000000000000",
19918 => "000000000000000000000000",
19919 => "000000000000000000000000",
19920 => "000000000000000000000000",
19921 => "000000000000000000000000",
19922 => "000000000000000000000000",
19923 => "000000000000000000000000",
19924 => "000000000000000000000000",
19925 => "000000000000000000000000",
19926 => "000000000000000000000000",
19927 => "000000000000000000000000",
19928 => "000000000000000000000000",
19929 => "000000000000000000000000",
19930 => "000000000000000000000000",
19931 => "000000000000000000000000",
19932 => "000000000000000000000000",
19933 => "000000000000000000000000",
19934 => "000000000000000000000000",
19935 => "000000000000000000000000",
19936 => "000000000000000000000000",
19937 => "000000000000000000000000",
19938 => "000000000000000000000000",
19939 => "000000000000000000000000",
19940 => "000000000000000000000000",
19941 => "000000000000000000000000",
19942 => "000000000000000000000000",
19943 => "000000000000000000000000",
19944 => "000000000000000000000000",
19945 => "000000000000000000000000",
19946 => "000000000000000000000000",
19947 => "000000000000000000000000",
19948 => "000000000000000000000000",
19949 => "000000000000000000000000",
19950 => "000000000000000000000000",
19951 => "000000000000000000000000",
19952 => "000000000000000000000000",
19953 => "000000000000000000000000",
19954 => "000000000000000000000000",
19955 => "000000000000000000000000",
19956 => "000000000000000000000000",
19957 => "000000000000000000000000",
19958 => "000000000000000000000000",
19959 => "000000000000000000000000",
19960 => "000000000000000000000000",
19961 => "000000000000000000000000",
19962 => "000000000000000000000000",
19963 => "000000000000000000000000",
19964 => "000000000000000000000000",
19965 => "000000000000000000000000",
19966 => "000000000000000000000000",
19967 => "000000000000000000000000",
19968 => "000000000000000000000000",
19969 => "000000000000000000000000",
19970 => "000000000000000000000000",
19971 => "000000000000000000000000",
19972 => "000000000000000000000000",
19973 => "000000000000000000000000",
19974 => "000000000000000000000000",
19975 => "000000000000000000000000",
19976 => "000000000000000000000000",
19977 => "000000000000000000000000",
19978 => "000000000000000000000000",
19979 => "000000000000000000000000",
19980 => "000000000000000000000000",
19981 => "000000000000000000000000",
19982 => "000000000000000000000000",
19983 => "000000000000000000000000",
19984 => "000000000000000000000000",
19985 => "000110010001100100011001",
19986 => "000110110001101100011011",
19987 => "001011110010111100101111",
19988 => "010000110100001101000011",
19989 => "010010000100100001001000",
19990 => "011001100110011001100110",
19991 => "011001100110011001100110",
19992 => "010001110100011101000111",
19993 => "010000110100001101000011",
19994 => "010000110100001101000011",
19995 => "010000110100001101000011",
19996 => "010000110100001101000011",
19997 => "010000110100001101000011",
19998 => "010000110100001101000011",
19999 => "010000110100001101000011",
20000 => "010000110100001101000011",
20001 => "001101110011011100110111",
20002 => "001010000010100000101000",
20003 => "001001000010010000100100",
20004 => "000000000000000000000000",
20005 => "000000000000000000000000",
20006 => "000000000000000000000000",
20007 => "000000000000000000000000",
20008 => "000000000000000000000000",
20009 => "000000000000000000000000",
20010 => "000001110000011000000100",
20011 => "011100000110010000111101",
20012 => "011100000110010000111101",
20013 => "011100000110010000111101",
20014 => "011100000110010000111101",
20015 => "010001100011111000100110",
20016 => "000000000000000000000000",
20017 => "000000000000000000000000",
20018 => "000000000000000000000000",
20019 => "000000000000000000000000",
20020 => "000000000000000000000000",
20021 => "000000000000000000000000",
20022 => "001001110010001000010101",
20023 => "011100000110010000111101",
20024 => "011100000110010000111101",
20025 => "011100000110010000111101",
20026 => "011100000110010000111101",
20027 => "001001110010001000010101",
20028 => "000000000000000000000000",
20029 => "000000000000000000000000",
20030 => "000000000000000000000000",
20031 => "000000000000000000000000",
20032 => "000000000000000000000000",
20033 => "000000000000000000000000",
20034 => "000110010001100100011001",
20035 => "001010000010100000101000",
20036 => "001011110010111100101111",
20037 => "010000110100001101000011",
20038 => "010000110100001101000011",
20039 => "010000110100001101000011",
20040 => "010000110100001101000011",
20041 => "010000110100001101000011",
20042 => "010000110100001101000011",
20043 => "010011000100110001001100",
20044 => "011001100110011001100110",
20045 => "011001100110011001100110",
20046 => "010001000100010001000100",
20047 => "010000110100001101000011",
20048 => "010000110100001101000011",
20049 => "010000110100001101000011",
20050 => "001110100011101000111010",
20051 => "000110110001101100011011",
20052 => "000110110001101100011011",
20053 => "000000010000000100000001",
20054 => "000000000000000000000000",
20055 => "000000000000000000000000",
20056 => "000000000000000000000000",
20057 => "000000000000000000000000",
20058 => "000000000000000000000000",
20059 => "000000000000000000000000",
20060 => "000000000000000000000000",
20061 => "000000000000000000000000",
20062 => "000000000000000000000000",
20063 => "000000000000000000000000",
20064 => "000000000000000000000000",
20065 => "000000000000000000000000",
20066 => "000000000000000000000000",
20067 => "000000000000000000000000",
20068 => "000000000000000000000000",
20069 => "000000000000000000000000",
20070 => "000000000000000000000000",
20071 => "000000000000000000000000",
20072 => "000000000000000000000000",
20073 => "000000000000000000000000",
20074 => "000000000000000000000000",
20075 => "000000000000000000000000",
20076 => "000000000000000000000000",
20077 => "000000000000000000000000",
20078 => "000000000000000000000000",
20079 => "000000000000000000000000",
20080 => "000000000000000000000000",
20081 => "000000000000000000000000",
20082 => "000000000000000000000000",
20083 => "000000000000000000000000",
20084 => "000000000000000000000000",
20085 => "000000000000000000000000",
20086 => "000000000000000000000000",
20087 => "000000000000000000000000",
20088 => "000000000000000000000000",
20089 => "000000000000000000000000",
20090 => "000000000000000000000000",
20091 => "000000000000000000000000",
20092 => "000000000000000000000000",
20093 => "000000000000000000000000",
20094 => "000000000000000000000000",
20095 => "000000000000000000000000",
20096 => "000000000000000000000000",
20097 => "000000000000000000000000",
20098 => "000000000000000000000000",
20099 => "000000000000000000000000",
20100 => "000000000000000000000000",
20101 => "000000000000000000000000",
20102 => "000000000000000000000000",
20103 => "000000000000000000000000",
20104 => "000000000000000000000000",
20105 => "000000000000000000000000",
20106 => "000000000000000000000000",
20107 => "000000000000000000000000",
20108 => "000000000000000000000000",
20109 => "000000000000000000000000",
20110 => "000000000000000000000000",
20111 => "000000000000000000000000",
20112 => "000000000000000000000000",
20113 => "000000000000000000000000",
20114 => "000000000000000000000000",
20115 => "000000000000000000000000",
20116 => "000000000000000000000000",
20117 => "000000000000000000000000",
20118 => "000000000000000000000000",
20119 => "000000000000000000000000",
20120 => "000000000000000000000000",
20121 => "000000000000000000000000",
20122 => "000000000000000000000000",
20123 => "000000000000000000000000",
20124 => "000000000000000000000000",
20125 => "000000000000000000000000",
20126 => "000000000000000000000000",
20127 => "000000000000000000000000",
20128 => "000000000000000000000000",
20129 => "000000000000000000000000",
20130 => "000000000000000000000000",
20131 => "000000000000000000000000",
20132 => "000000000000000000000000",
20133 => "000000000000000000000000",
20134 => "000000000000000000000000",
20135 => "001111010011110100111101",
20136 => "010000110100001101000011",
20137 => "010000110100001101000011",
20138 => "010000110100001101000011",
20139 => "010010000100100001001000",
20140 => "011001100110011001100110",
20141 => "011001100110011001100110",
20142 => "010001110100011101000111",
20143 => "010000110100001101000011",
20144 => "010000110100001101000011",
20145 => "010000110100001101000011",
20146 => "010000110100001101000011",
20147 => "010000110100001101000011",
20148 => "010000110100001101000011",
20149 => "010000110100001101000011",
20150 => "010000110100001101000011",
20151 => "001001100010011000100110",
20152 => "000000000000000000000000",
20153 => "000000000000000000000000",
20154 => "000000000000000000000000",
20155 => "000000000000000000000000",
20156 => "000000000000000000000000",
20157 => "000000000000000000000000",
20158 => "000000000000000000000000",
20159 => "000000000000000000000000",
20160 => "000010000000011000000000",
20161 => "011111110110000000000000",
20162 => "011111110110000000000000",
20163 => "011111110110000000000000",
20164 => "011111110110000000000000",
20165 => "010011110011110000000000",
20166 => "000000000000000000000000",
20167 => "000000000000000000000000",
20168 => "000000000000000000000000",
20169 => "000000000000000000000000",
20170 => "000000000000000000000000",
20171 => "000000000000000000000000",
20172 => "001011000010000100000000",
20173 => "011111110110000000000000",
20174 => "011111110110000000000000",
20175 => "011111110110000000000000",
20176 => "011111110110000000000000",
20177 => "001011000010000100000000",
20178 => "000000000000000000000000",
20179 => "000000000000000000000000",
20180 => "000000000000000000000000",
20181 => "000000000000000000000000",
20182 => "000000000000000000000000",
20183 => "000000000000000000000000",
20184 => "000000000000000000000000",
20185 => "000000000000000000000000",
20186 => "000100110001001100010011",
20187 => "010000110100001101000011",
20188 => "010000110100001101000011",
20189 => "010000110100001101000011",
20190 => "010000110100001101000011",
20191 => "010000110100001101000011",
20192 => "010000110100001101000011",
20193 => "010011000100110001001100",
20194 => "011001100110011001100110",
20195 => "011001100110011001100110",
20196 => "010001000100010001000100",
20197 => "010000110100001101000011",
20198 => "010000110100001101000011",
20199 => "010000110100001101000011",
20200 => "010000110100001101000011",
20201 => "010000110100001101000011",
20202 => "010000110100001101000011",
20203 => "000001000000010000000100",
20204 => "000000000000000000000000",
20205 => "000000000000000000000000",
20206 => "000000000000000000000000",
20207 => "000000000000000000000000",
20208 => "000000000000000000000000",
20209 => "000000000000000000000000",
20210 => "000000000000000000000000",
20211 => "000000000000000000000000",
20212 => "000000000000000000000000",
20213 => "000000000000000000000000",
20214 => "000000000000000000000000",
20215 => "000000000000000000000000",
20216 => "000000000000000000000000",
20217 => "000000000000000000000000",
20218 => "000000000000000000000000",
20219 => "000000000000000000000000",
20220 => "000000000000000000000000",
20221 => "000000000000000000000000",
20222 => "000000000000000000000000",
20223 => "000000000000000000000000",
20224 => "000000000000000000000000",
20225 => "000000000000000000000000",
20226 => "000000000000000000000000",
20227 => "000000000000000000000000",
20228 => "000000000000000000000000",
20229 => "000000000000000000000000",
20230 => "000000000000000000000000",
20231 => "000000000000000000000000",
20232 => "000000000000000000000000",
20233 => "000000000000000000000000",
20234 => "000000000000000000000000",
20235 => "000000000000000000000000",
20236 => "000000000000000000000000",
20237 => "000000000000000000000000",
20238 => "000000000000000000000000",
20239 => "000000000000000000000000",
20240 => "000000000000000000000000",
20241 => "000000000000000000000000",
20242 => "000000000000000000000000",
20243 => "000000000000000000000000",
20244 => "000000000000000000000000",
20245 => "000000000000000000000000",
20246 => "000000000000000000000000",
20247 => "000000000000000000000000",
20248 => "000000000000000000000000",
20249 => "000000000000000000000000",
20250 => "000000000000000000000000",
20251 => "000000000000000000000000",
20252 => "000000000000000000000000",
20253 => "000000000000000000000000",
20254 => "000000000000000000000000",
20255 => "000000000000000000000000",
20256 => "000000000000000000000000",
20257 => "000000000000000000000000",
20258 => "000000000000000000000000",
20259 => "000000000000000000000000",
20260 => "000000000000000000000000",
20261 => "000000000000000000000000",
20262 => "000000000000000000000000",
20263 => "000000000000000000000000",
20264 => "000000000000000000000000",
20265 => "000000000000000000000000",
20266 => "000000000000000000000000",
20267 => "000000000000000000000000",
20268 => "000000000000000000000000",
20269 => "000000000000000000000000",
20270 => "000000000000000000000000",
20271 => "000000000000000000000000",
20272 => "000000000000000000000000",
20273 => "000000000000000000000000",
20274 => "000000000000000000000000",
20275 => "000000000000000000000000",
20276 => "000000000000000000000000",
20277 => "000000000000000000000000",
20278 => "000000000000000000000000",
20279 => "000000000000000000000000",
20280 => "000000000000000000000000",
20281 => "000000000000000000000000",
20282 => "000000010000000100000001",
20283 => "000001000000010000000100",
20284 => "000001000000010000000100",
20285 => "001111100011111000111110",
20286 => "010000110100001101000011",
20287 => "010000110100001101000011",
20288 => "010000110100001101000011",
20289 => "010010000100100001001000",
20290 => "011001100110011001100110",
20291 => "011001100110011001100110",
20292 => "010001110100011101000111",
20293 => "010000110100001101000011",
20294 => "010000110100001101000011",
20295 => "010000110100001101000011",
20296 => "010000110100001101000011",
20297 => "010000110100001101000011",
20298 => "010000110100001101000011",
20299 => "010000110100001101000011",
20300 => "010000110100001101000011",
20301 => "001001100010011000100110",
20302 => "000000000000000000000000",
20303 => "000000000000000000000000",
20304 => "000000000000000000000000",
20305 => "000000000000000000000000",
20306 => "000000000000000000000000",
20307 => "000000000000000000000000",
20308 => "000000000000000000000000",
20309 => "000000000000000000000000",
20310 => "000001110000011000000000",
20311 => "011101110101101000000000",
20312 => "011101110101101000000000",
20313 => "011101110101101000000000",
20314 => "011101110101101000000000",
20315 => "010010100011100000000000",
20316 => "000000000000000000000000",
20317 => "000000000000000000000000",
20318 => "000000000000000000000000",
20319 => "000000000000000000000000",
20320 => "000000000000000000000000",
20321 => "000000000000000000000000",
20322 => "001010010001111100000000",
20323 => "011101110101101000000000",
20324 => "011101110101101000000000",
20325 => "011101110101101000000000",
20326 => "011101110101101000000000",
20327 => "001010010001111100000000",
20328 => "000000000000000000000000",
20329 => "000000000000000000000000",
20330 => "000000000000000000000000",
20331 => "000000000000000000000000",
20332 => "000000000000000000000000",
20333 => "000000000000000000000000",
20334 => "000000000000000000000000",
20335 => "000000000000000000000000",
20336 => "000100110001001100010011",
20337 => "010000110100001101000011",
20338 => "010000110100001101000011",
20339 => "010000110100001101000011",
20340 => "010000110100001101000011",
20341 => "010000110100001101000011",
20342 => "010000110100001101000011",
20343 => "010011000100110001001100",
20344 => "011001100110011001100110",
20345 => "011001100110011001100110",
20346 => "010001000100010001000100",
20347 => "010000110100001101000011",
20348 => "010000110100001101000011",
20349 => "010000110100001101000011",
20350 => "010000110100001101000011",
20351 => "010000110100001101000011",
20352 => "010000110100001101000011",
20353 => "000010000000100000001000",
20354 => "000001000000010000000100",
20355 => "000000100000001000000010",
20356 => "000000000000000000000000",
20357 => "000000000000000000000000",
20358 => "000000000000000000000000",
20359 => "000000000000000000000000",
20360 => "000000000000000000000000",
20361 => "000000000000000000000000",
20362 => "000000000000000000000000",
20363 => "000000000000000000000000",
20364 => "000000000000000000000000",
20365 => "000000000000000000000000",
20366 => "000000000000000000000000",
20367 => "000000000000000000000000",
20368 => "000000000000000000000000",
20369 => "000000000000000000000000",
20370 => "000000000000000000000000",
20371 => "000000000000000000000000",
20372 => "000000000000000000000000",
20373 => "000000000000000000000000",
20374 => "000000000000000000000000",
20375 => "000000000000000000000000",
20376 => "000000000000000000000000",
20377 => "000000000000000000000000",
20378 => "000000000000000000000000",
20379 => "000000000000000000000000",
20380 => "000000000000000000000000",
20381 => "000000000000000000000000",
20382 => "000000000000000000000000",
20383 => "000000000000000000000000",
20384 => "000000000000000000000000",
20385 => "000000000000000000000000",
20386 => "000000000000000000000000",
20387 => "000000000000000000000000",
20388 => "000000000000000000000000",
20389 => "000000000000000000000000",
20390 => "000000000000000000000000",
20391 => "000000000000000000000000",
20392 => "000000000000000000000000",
20393 => "000000000000000000000000",
20394 => "000000000000000000000000",
20395 => "000000000000000000000000",
20396 => "000000000000000000000000",
20397 => "000000000000000000000000",
20398 => "000000000000000000000000",
20399 => "000000000000000000000000",
20400 => "000000000000000000000000",
20401 => "000000000000000000000000",
20402 => "000000000000000000000000",
20403 => "000000000000000000000000",
20404 => "000000000000000000000000",
20405 => "000000000000000000000000",
20406 => "000000000000000000000000",
20407 => "000000000000000000000000",
20408 => "000000000000000000000000",
20409 => "000000000000000000000000",
20410 => "000000000000000000000000",
20411 => "000000000000000000000000",
20412 => "000000000000000000000000",
20413 => "000000000000000000000000",
20414 => "000000000000000000000000",
20415 => "000000000000000000000000",
20416 => "000000000000000000000000",
20417 => "000000000000000000000000",
20418 => "000000000000000000000000",
20419 => "000000000000000000000000",
20420 => "000000000000000000000000",
20421 => "000000000000000000000000",
20422 => "000000000000000000000000",
20423 => "000000000000000000000000",
20424 => "000000000000000000000000",
20425 => "000000000000000000000000",
20426 => "000000000000000000000000",
20427 => "000000000000000000000000",
20428 => "000000000000000000000000",
20429 => "000000000000000000000000",
20430 => "000000000000000000000000",
20431 => "000000000000000000000000",
20432 => "000011010000110100001101",
20433 => "010000110100001101000011",
20434 => "010000110100001101000011",
20435 => "010000110100001101000011",
20436 => "010000110100001101000011",
20437 => "010000110100001101000011",
20438 => "010000110100001101000011",
20439 => "010010000100100001001000",
20440 => "011001100110011001100110",
20441 => "011001100110011001100110",
20442 => "010001110100011101000111",
20443 => "010000110100001101000011",
20444 => "010000110100001101000011",
20445 => "010000110100001101000011",
20446 => "010000110100001101000011",
20447 => "010000110100001101000011",
20448 => "010000110100001101000011",
20449 => "010000110100001101000011",
20450 => "010000110100001101000011",
20451 => "001001100010011000100110",
20452 => "000000000000000000000000",
20453 => "000000000000000000000000",
20454 => "000000000000000000000000",
20455 => "000000000000000000000000",
20456 => "000000000000000000000000",
20457 => "000000000000000000000000",
20458 => "000000000000000000000000",
20459 => "000000000000000000000000",
20460 => "000000000000000000000000",
20461 => "000000000000000000000000",
20462 => "000000000000000000000000",
20463 => "000000000000000000000000",
20464 => "000000000000000000000000",
20465 => "000000000000000000000000",
20466 => "000000000000000000000000",
20467 => "000000000000000000000000",
20468 => "000000000000000000000000",
20469 => "000000000000000000000000",
20470 => "000000000000000000000000",
20471 => "000000000000000000000000",
20472 => "000000000000000000000000",
20473 => "000000000000000000000000",
20474 => "000000000000000000000000",
20475 => "000000000000000000000000",
20476 => "000000000000000000000000",
20477 => "000000000000000000000000",
20478 => "000000000000000000000000",
20479 => "000000000000000000000000",
20480 => "000000000000000000000000",
20481 => "000000000000000000000000",
20482 => "000000000000000000000000",
20483 => "000000000000000000000000",
20484 => "000000000000000000000000",
20485 => "000000000000000000000000",
20486 => "000100110001001100010011",
20487 => "010000110100001101000011",
20488 => "010000110100001101000011",
20489 => "010000110100001101000011",
20490 => "010000110100001101000011",
20491 => "010000110100001101000011",
20492 => "010000110100001101000011",
20493 => "010011000100110001001100",
20494 => "011001100110011001100110",
20495 => "011001100110011001100110",
20496 => "010001000100010001000100",
20497 => "010000110100001101000011",
20498 => "010000110100001101000011",
20499 => "010000110100001101000011",
20500 => "010000110100001101000011",
20501 => "010000110100001101000011",
20502 => "010000110100001101000011",
20503 => "010000110100001101000011",
20504 => "010000110100001101000011",
20505 => "000111110001111100011111",
20506 => "000000000000000000000000",
20507 => "000000000000000000000000",
20508 => "000000000000000000000000",
20509 => "000000000000000000000000",
20510 => "000000000000000000000000",
20511 => "000000000000000000000000",
20512 => "000000000000000000000000",
20513 => "000000000000000000000000",
20514 => "000000000000000000000000",
20515 => "000000000000000000000000",
20516 => "000000000000000000000000",
20517 => "000000000000000000000000",
20518 => "000000000000000000000000",
20519 => "000000000000000000000000",
20520 => "000000000000000000000000",
20521 => "000000000000000000000000",
20522 => "000000000000000000000000",
20523 => "000000000000000000000000",
20524 => "000000000000000000000000",
20525 => "000000000000000000000000",
20526 => "000000000000000000000000",
20527 => "000000000000000000000000",
20528 => "000000000000000000000000",
20529 => "000000000000000000000000",
20530 => "000000000000000000000000",
20531 => "000000000000000000000000",
20532 => "000000000000000000000000",
20533 => "000000000000000000000000",
20534 => "000000000000000000000000",
20535 => "000000000000000000000000",
20536 => "000000000000000000000000",
20537 => "000000000000000000000000",
20538 => "000000000000000000000000",
20539 => "000000000000000000000000",
20540 => "000000000000000000000000",
20541 => "000000000000000000000000",
20542 => "000000000000000000000000",
20543 => "000000000000000000000000",
20544 => "000000000000000000000000",
20545 => "000000000000000000000000",
20546 => "000000000000000000000000",
20547 => "000000000000000000000000",
20548 => "000000000000000000000000",
20549 => "000000000000000000000000",
20550 => "000000000000000000000000",
20551 => "000000000000000000000000",
20552 => "000000000000000000000000",
20553 => "000000000000000000000000",
20554 => "000000000000000000000000",
20555 => "000000000000000000000000",
20556 => "000000000000000000000000",
20557 => "000000000000000000000000",
20558 => "000000000000000000000000",
20559 => "000000000000000000000000",
20560 => "000000000000000000000000",
20561 => "000000000000000000000000",
20562 => "000000000000000000000000",
20563 => "000000000000000000000000",
20564 => "000000000000000000000000",
20565 => "000000000000000000000000",
20566 => "000000000000000000000000",
20567 => "000000000000000000000000",
20568 => "000000000000000000000000",
20569 => "000000000000000000000000",
20570 => "000000000000000000000000",
20571 => "000000000000000000000000",
20572 => "000000000000000000000000",
20573 => "000000000000000000000000",
20574 => "000000000000000000000000",
20575 => "000000000000000000000000",
20576 => "000000000000000000000000",
20577 => "000000000000000000000000",
20578 => "000000000000000000000000",
20579 => "000000000000000000000000",
20580 => "000000000000000000000000",
20581 => "000000000000000000000000",
20582 => "000011010000110100001101",
20583 => "010000110100001101000011",
20584 => "010000110100001101000011",
20585 => "010000110100001101000011",
20586 => "010000110100001101000011",
20587 => "010000110100001101000011",
20588 => "010000110100001101000011",
20589 => "010010000100100001001000",
20590 => "011001100110011001100110",
20591 => "011001100110011001100110",
20592 => "010001110100011101000111",
20593 => "010000110100001101000011",
20594 => "010000110100001101000011",
20595 => "010000110100001101000011",
20596 => "010000110100001101000011",
20597 => "010000110100001101000011",
20598 => "010000110100001101000011",
20599 => "010000110100001101000011",
20600 => "010000110100001101000011",
20601 => "001001100010011000100110",
20602 => "000000000000000000000000",
20603 => "000000000000000000000000",
20604 => "000000000000000000000000",
20605 => "000000000000000000000000",
20606 => "000000000000000000000000",
20607 => "000000000000000000000000",
20608 => "000000000000000000000000",
20609 => "000000000000000000000000",
20610 => "000000000000000000000000",
20611 => "000000000000000000000000",
20612 => "000000000000000000000000",
20613 => "000000000000000000000000",
20614 => "000000000000000000000000",
20615 => "000000000000000000000000",
20616 => "000000000000000000000000",
20617 => "000000000000000000000000",
20618 => "000000000000000000000000",
20619 => "000000000000000000000000",
20620 => "000000000000000000000000",
20621 => "000000000000000000000000",
20622 => "000000000000000000000000",
20623 => "000000000000000000000000",
20624 => "000000000000000000000000",
20625 => "000000000000000000000000",
20626 => "000000000000000000000000",
20627 => "000000000000000000000000",
20628 => "000000000000000000000000",
20629 => "000000000000000000000000",
20630 => "000000000000000000000000",
20631 => "000000000000000000000000",
20632 => "000000000000000000000000",
20633 => "000000000000000000000000",
20634 => "000000000000000000000000",
20635 => "000000000000000000000000",
20636 => "000100110001001100010011",
20637 => "010000110100001101000011",
20638 => "010000110100001101000011",
20639 => "010000110100001101000011",
20640 => "010000110100001101000011",
20641 => "010000110100001101000011",
20642 => "010000110100001101000011",
20643 => "010011000100110001001100",
20644 => "011001100110011001100110",
20645 => "011001100110011001100110",
20646 => "010001000100010001000100",
20647 => "010000110100001101000011",
20648 => "010000110100001101000011",
20649 => "010000110100001101000011",
20650 => "010000110100001101000011",
20651 => "010000110100001101000011",
20652 => "010000110100001101000011",
20653 => "010000110100001101000011",
20654 => "010000110100001101000011",
20655 => "000111110001111100011111",
20656 => "000000000000000000000000",
20657 => "000000000000000000000000",
20658 => "000000000000000000000000",
20659 => "000000000000000000000000",
20660 => "000000000000000000000000",
20661 => "000000000000000000000000",
20662 => "000000000000000000000000",
20663 => "000000000000000000000000",
20664 => "000000000000000000000000",
20665 => "000000000000000000000000",
20666 => "000000000000000000000000",
20667 => "000000000000000000000000",
20668 => "000000000000000000000000",
20669 => "000000000000000000000000",
20670 => "000000000000000000000000",
20671 => "000000000000000000000000",
20672 => "000000000000000000000000",
20673 => "000000000000000000000000",
20674 => "000000000000000000000000",
20675 => "000000000000000000000000",
20676 => "000000000000000000000000",
20677 => "000000000000000000000000",
20678 => "000000000000000000000000",
20679 => "000000000000000000000000",
20680 => "000000000000000000000000",
20681 => "000000000000000000000000",
20682 => "000000000000000000000000",
20683 => "000000000000000000000000",
20684 => "000000000000000000000000",
20685 => "000000000000000000000000",
20686 => "000000000000000000000000",
20687 => "000000000000000000000000",
20688 => "000000000000000000000000",
20689 => "000000000000000000000000",
20690 => "000000000000000000000000",
20691 => "000000000000000000000000",
20692 => "000000000000000000000000",
20693 => "000000000000000000000000",
20694 => "000000000000000000000000",
20695 => "000000000000000000000000",
20696 => "000000000000000000000000",
20697 => "000000000000000000000000",
20698 => "000000000000000000000000",
20699 => "000000000000000000000000",
20700 => "000000000000000000000000",
20701 => "000000000000000000000000",
20702 => "000000000000000000000000",
20703 => "000000000000000000000000",
20704 => "000000000000000000000000",
20705 => "000000000000000000000000",
20706 => "000000000000000000000000",
20707 => "000000000000000000000000",
20708 => "000000000000000000000000",
20709 => "000000000000000000000000",
20710 => "000000000000000000000000",
20711 => "000000000000000000000000",
20712 => "000000000000000000000000",
20713 => "000000000000000000000000",
20714 => "000000000000000000000000",
20715 => "000000000000000000000000",
20716 => "000000000000000000000000",
20717 => "000000000000000000000000",
20718 => "000000000000000000000000",
20719 => "000000000000000000000000",
20720 => "000000000000000000000000",
20721 => "000000000000000000000000",
20722 => "000000000000000000000000",
20723 => "000000000000000000000000",
20724 => "000000000000000000000000",
20725 => "000000000000000000000000",
20726 => "000000000000000000000000",
20727 => "000000000000000000000000",
20728 => "000000000000000000000000",
20729 => "000000000000000000000000",
20730 => "000110100001101000011010",
20731 => "001100010011000100110001",
20732 => "001101000011010000110100",
20733 => "010000110100001101000011",
20734 => "010000110100001101000011",
20735 => "010000110100001101000011",
20736 => "010000110100001101000011",
20737 => "010000110100001101000011",
20738 => "010000110100001101000011",
20739 => "010001000100010001000100",
20740 => "010011000100110001001100",
20741 => "010011000100110001001100",
20742 => "010001000100010001000100",
20743 => "010000110100001101000011",
20744 => "010000110100001101000011",
20745 => "010000110100001101000011",
20746 => "010000110100001101000011",
20747 => "010000110100001101000011",
20748 => "010000110100001101000011",
20749 => "000110100001101000011010",
20750 => "000100100001001000010010",
20751 => "000010100000101000001010",
20752 => "000000000000000000000000",
20753 => "000000000000000000000000",
20754 => "000000000000000000000000",
20755 => "000000000000000000000000",
20756 => "000000000000000000000000",
20757 => "000000000000000000000000",
20758 => "000000000000000000000000",
20759 => "000000000000000000000000",
20760 => "000010110000100000000101",
20761 => "101101001000001001001110",
20762 => "101101001000001001001110",
20763 => "101110001010101100010101",
20764 => "101110101011101000000000",
20765 => "011101000111010000000000",
20766 => "000000000000000000000000",
20767 => "000000000000000000000000",
20768 => "000000000000000000000000",
20769 => "000000000000000000000000",
20770 => "000000000000000000000000",
20771 => "000000000000000000000000",
20772 => "010000000100000000000000",
20773 => "101110101011101000000000",
20774 => "101110101011101000000000",
20775 => "101101001000001001001110",
20776 => "101101001000001001001110",
20777 => "001111100010110100011011",
20778 => "000000000000000000000000",
20779 => "000000000000000000000000",
20780 => "000000000000000000000000",
20781 => "000000000000000000000000",
20782 => "000000000000000000000000",
20783 => "000000000000000000000000",
20784 => "000000000000000000000000",
20785 => "000000000000000000000000",
20786 => "000001010000010100000101",
20787 => "000100100001001000010010",
20788 => "000100100001001000010010",
20789 => "010000100100001001000010",
20790 => "010000110100001101000011",
20791 => "010000110100001101000011",
20792 => "010000110100001101000011",
20793 => "010001010100010101000101",
20794 => "010011000100110001001100",
20795 => "010011000100110001001100",
20796 => "010000110100001101000011",
20797 => "010000110100001101000011",
20798 => "010000110100001101000011",
20799 => "010000110100001101000011",
20800 => "010000110100001101000011",
20801 => "010000110100001101000011",
20802 => "010000110100001101000011",
20803 => "010000110100001101000011",
20804 => "010000110100001101000011",
20805 => "001110010011100100111001",
20806 => "001100010011000100110001",
20807 => "001010000010100000101000",
20808 => "000000000000000000000000",
20809 => "000000000000000000000000",
20810 => "000000000000000000000000",
20811 => "000000000000000000000000",
20812 => "000000000000000000000000",
20813 => "000000000000000000000000",
20814 => "000000000000000000000000",
20815 => "000000000000000000000000",
20816 => "000000000000000000000000",
20817 => "000000000000000000000000",
20818 => "000000000000000000000000",
20819 => "000000000000000000000000",
20820 => "000000000000000000000000",
20821 => "000000000000000000000000",
20822 => "000000000000000000000000",
20823 => "000000000000000000000000",
20824 => "000000000000000000000000",
20825 => "000000000000000000000000",
20826 => "000000000000000000000000",
20827 => "000000000000000000000000",
20828 => "000000000000000000000000",
20829 => "000000000000000000000000",
20830 => "000000000000000000000000",
20831 => "000000000000000000000000",
20832 => "000000000000000000000000",
20833 => "000000000000000000000000",
20834 => "000000000000000000000000",
20835 => "000000000000000000000000",
20836 => "000000000000000000000000",
20837 => "000000000000000000000000",
20838 => "000000000000000000000000",
20839 => "000000000000000000000000",
20840 => "000000000000000000000000",
20841 => "000000000000000000000000",
20842 => "000000000000000000000000",
20843 => "000000000000000000000000",
20844 => "000000000000000000000000",
20845 => "000000000000000000000000",
20846 => "000000000000000000000000",
20847 => "000000000000000000000000",
20848 => "000000000000000000000000",
20849 => "000000000000000000000000",
20850 => "000000000000000000000000",
20851 => "000000000000000000000000",
20852 => "000000000000000000000000",
20853 => "000000000000000000000000",
20854 => "000000000000000000000000",
20855 => "000000000000000000000000",
20856 => "000000000000000000000000",
20857 => "000000000000000000000000",
20858 => "000000000000000000000000",
20859 => "000000000000000000000000",
20860 => "000000000000000000000000",
20861 => "000000000000000000000000",
20862 => "000000000000000000000000",
20863 => "000000000000000000000000",
20864 => "000000000000000000000000",
20865 => "000000000000000000000000",
20866 => "000000000000000000000000",
20867 => "000000000000000000000000",
20868 => "000000000000000000000000",
20869 => "000000000000000000000000",
20870 => "000000000000000000000000",
20871 => "000000000000000000000000",
20872 => "000000000000000000000000",
20873 => "000000000000000000000000",
20874 => "000000000000000000000000",
20875 => "000000000000000000000000",
20876 => "000000000000000000000000",
20877 => "000000000000000000000000",
20878 => "000000000000000000000000",
20879 => "000000000000000000000000",
20880 => "001001000010010000100100",
20881 => "010000110100001101000011",
20882 => "010000110100001101000011",
20883 => "010000110100001101000011",
20884 => "010000110100001101000011",
20885 => "010000110100001101000011",
20886 => "010000110100001101000011",
20887 => "010000110100001101000011",
20888 => "010000110100001101000011",
20889 => "010000110100001101000011",
20890 => "010000110100001101000011",
20891 => "010000110100001101000011",
20892 => "010000110100001101000011",
20893 => "010000110100001101000011",
20894 => "010000110100001101000011",
20895 => "010000110100001101000011",
20896 => "010000110100001101000011",
20897 => "010000110100001101000011",
20898 => "010000110100001101000011",
20899 => "000010110000101100001011",
20900 => "000000000000000000000000",
20901 => "000000000000000000000000",
20902 => "000000000000000000000000",
20903 => "000000000000000000000000",
20904 => "000000000000000000000000",
20905 => "000000000000000000000000",
20906 => "000000000000000000000000",
20907 => "000000000000000000000000",
20908 => "000000000000000000000000",
20909 => "000000000000000000000000",
20910 => "000011110000101100000111",
20911 => "111101101011001001101011",
20912 => "111101101011001001101011",
20913 => "111111011110101000011101",
20914 => "111111111111111100000000",
20915 => "100111111001111100000000",
20916 => "000000000000000000000000",
20917 => "000000000000000000000000",
20918 => "000000000000000000000000",
20919 => "000000000000000000000000",
20920 => "000000000000000000000000",
20921 => "000000000000000000000000",
20922 => "010110000101100000000000",
20923 => "111111111111111100000000",
20924 => "111111111111111100000000",
20925 => "111101101011001001101011",
20926 => "111101101011001001101011",
20927 => "010101010011110100100101",
20928 => "000000000000000000000000",
20929 => "000000000000000000000000",
20930 => "000000000000000000000000",
20931 => "000000000000000000000000",
20932 => "000000000000000000000000",
20933 => "000000000000000000000000",
20934 => "000000000000000000000000",
20935 => "000000000000000000000000",
20936 => "000000000000000000000000",
20937 => "000000000000000000000000",
20938 => "000000000000000000000000",
20939 => "010000100100001001000010",
20940 => "010000110100001101000011",
20941 => "010000110100001101000011",
20942 => "010000110100001101000011",
20943 => "010000110100001101000011",
20944 => "010000110100001101000011",
20945 => "010000110100001101000011",
20946 => "010000110100001101000011",
20947 => "010000110100001101000011",
20948 => "010000110100001101000011",
20949 => "010000110100001101000011",
20950 => "010000110100001101000011",
20951 => "010000110100001101000011",
20952 => "010000110100001101000011",
20953 => "010000110100001101000011",
20954 => "010000110100001101000011",
20955 => "010000110100001101000011",
20956 => "010000110100001101000011",
20957 => "001101100011011000110110",
20958 => "000000000000000000000000",
20959 => "000000000000000000000000",
20960 => "000000000000000000000000",
20961 => "000000000000000000000000",
20962 => "000000000000000000000000",
20963 => "000000000000000000000000",
20964 => "000000000000000000000000",
20965 => "000000000000000000000000",
20966 => "000000000000000000000000",
20967 => "000000000000000000000000",
20968 => "000000000000000000000000",
20969 => "000000000000000000000000",
20970 => "000000000000000000000000",
20971 => "000000000000000000000000",
20972 => "000000000000000000000000",
20973 => "000000000000000000000000",
20974 => "000000000000000000000000",
20975 => "000000000000000000000000",
20976 => "000000000000000000000000",
20977 => "000000000000000000000000",
20978 => "000000000000000000000000",
20979 => "000000000000000000000000",
20980 => "000000000000000000000000",
20981 => "000000000000000000000000",
20982 => "000000000000000000000000",
20983 => "000000000000000000000000",
20984 => "000000000000000000000000",
20985 => "000000000000000000000000",
20986 => "000000000000000000000000",
20987 => "000000000000000000000000",
20988 => "000000000000000000000000",
20989 => "000000000000000000000000",
20990 => "000000000000000000000000",
20991 => "000000000000000000000000",
20992 => "000000000000000000000000",
20993 => "000000000000000000000000",
20994 => "000000000000000000000000",
20995 => "000000000000000000000000",
20996 => "000000000000000000000000",
20997 => "000000000000000000000000",
20998 => "000000000000000000000000",
20999 => "000000000000000000000000",
21000 => "000000000000000000000000",
21001 => "000000000000000000000000",
21002 => "000000000000000000000000",
21003 => "000000000000000000000000",
21004 => "000000000000000000000000",
21005 => "000000000000000000000000",
21006 => "000000000000000000000000",
21007 => "000000000000000000000000",
21008 => "000000000000000000000000",
21009 => "000000000000000000000000",
21010 => "000000000000000000000000",
21011 => "000000000000000000000000",
21012 => "000000000000000000000000",
21013 => "000000000000000000000000",
21014 => "000000000000000000000000",
21015 => "000000000000000000000000",
21016 => "000000000000000000000000",
21017 => "000000000000000000000000",
21018 => "000000000000000000000000",
21019 => "000000000000000000000000",
21020 => "000000000000000000000000",
21021 => "000000000000000000000000",
21022 => "000000000000000000000000",
21023 => "000000000000000000000000",
21024 => "000000000000000000000000",
21025 => "000000000000000000000000",
21026 => "000000000000000000000000",
21027 => "000000000000000000000000",
21028 => "000000000000000000000000",
21029 => "000000000000000000000000",
21030 => "001001000010010000100100",
21031 => "010000110100001101000011",
21032 => "010000110100001101000011",
21033 => "010000110100001101000011",
21034 => "010000110100001101000011",
21035 => "010000110100001101000011",
21036 => "010000110100001101000011",
21037 => "010000110100001101000011",
21038 => "010000110100001101000011",
21039 => "010000110100001101000011",
21040 => "010000110100001101000011",
21041 => "010000110100001101000011",
21042 => "010000110100001101000011",
21043 => "010000110100001101000011",
21044 => "010000110100001101000011",
21045 => "010000110100001101000011",
21046 => "010000110100001101000011",
21047 => "010000110100001101000011",
21048 => "010000110100001101000011",
21049 => "000010110000101100001011",
21050 => "000000000000000000000000",
21051 => "000000000000000000000000",
21052 => "000000000000000000000000",
21053 => "000000000000000000000000",
21054 => "000000000000000000000000",
21055 => "000000000000000000000000",
21056 => "000000000000000000000000",
21057 => "000000000000000000000000",
21058 => "000000000000000000000000",
21059 => "000000000000000000000000",
21060 => "000011110000101100000111",
21061 => "111101101011001001101011",
21062 => "111101101011001001101011",
21063 => "111110101101010100111010",
21064 => "111111001110001000101000",
21065 => "100111011000110100011001",
21066 => "000000000000000000000000",
21067 => "000000000000000000000000",
21068 => "000000000000000000000000",
21069 => "000000000000000000000000",
21070 => "000000000000000000000000",
21071 => "000000000000000000000000",
21072 => "010101100100111000001110",
21073 => "111111001110001000101000",
21074 => "111111001110001000101000",
21075 => "100110100110111101000011",
21076 => "100110100110111101000011",
21077 => "001101010010011000010111",
21078 => "000000000000000000000000",
21079 => "000000000000000000000000",
21080 => "000000000000000000000000",
21081 => "000000000000000000000000",
21082 => "000000000000000000000000",
21083 => "000000000000000000000000",
21084 => "000000000000000000000000",
21085 => "000000000000000000000000",
21086 => "000000000000000000000000",
21087 => "000000000000000000000000",
21088 => "000000000000000000000000",
21089 => "010000100100001001000010",
21090 => "010000110100001101000011",
21091 => "010000110100001101000011",
21092 => "010000110100001101000011",
21093 => "010000110100001101000011",
21094 => "010000110100001101000011",
21095 => "010000110100001101000011",
21096 => "010000110100001101000011",
21097 => "010000110100001101000011",
21098 => "010000110100001101000011",
21099 => "010000110100001101000011",
21100 => "010000110100001101000011",
21101 => "010000110100001101000011",
21102 => "010000110100001101000011",
21103 => "010000110100001101000011",
21104 => "010000110100001101000011",
21105 => "010000110100001101000011",
21106 => "010000110100001101000011",
21107 => "001101100011011000110110",
21108 => "000000000000000000000000",
21109 => "000000000000000000000000",
21110 => "000000000000000000000000",
21111 => "000000000000000000000000",
21112 => "000000000000000000000000",
21113 => "000000000000000000000000",
21114 => "000000000000000000000000",
21115 => "000000000000000000000000",
21116 => "000000000000000000000000",
21117 => "000000000000000000000000",
21118 => "000000000000000000000000",
21119 => "000000000000000000000000",
21120 => "000000000000000000000000",
21121 => "000000000000000000000000",
21122 => "000000000000000000000000",
21123 => "000000000000000000000000",
21124 => "000000000000000000000000",
21125 => "000000000000000000000000",
21126 => "000000000000000000000000",
21127 => "000000000000000000000000",
21128 => "000000000000000000000000",
21129 => "000000000000000000000000",
21130 => "000000000000000000000000",
21131 => "000000000000000000000000",
21132 => "000000000000000000000000",
21133 => "000000000000000000000000",
21134 => "000000000000000000000000",
21135 => "000000000000000000000000",
21136 => "000000000000000000000000",
21137 => "000000000000000000000000",
21138 => "000000000000000000000000",
21139 => "000000000000000000000000",
21140 => "000000000000000000000000",
21141 => "000000000000000000000000",
21142 => "000000000000000000000000",
21143 => "000000000000000000000000",
21144 => "000000000000000000000000",
21145 => "000000000000000000000000",
21146 => "000000000000000000000000",
21147 => "000000000000000000000000",
21148 => "000000000000000000000000",
21149 => "000000000000000000000000",
21150 => "000000000000000000000000",
21151 => "000000000000000000000000",
21152 => "000000000000000000000000",
21153 => "000000000000000000000000",
21154 => "000000000000000000000000",
21155 => "000000000000000000000000",
21156 => "000000000000000000000000",
21157 => "000000000000000000000000",
21158 => "000000000000000000000000",
21159 => "000000000000000000000000",
21160 => "000000000000000000000000",
21161 => "000000000000000000000000",
21162 => "000000000000000000000000",
21163 => "000000000000000000000000",
21164 => "000000000000000000000000",
21165 => "000000000000000000000000",
21166 => "000000000000000000000000",
21167 => "000000000000000000000000",
21168 => "000000000000000000000000",
21169 => "000000000000000000000000",
21170 => "000000000000000000000000",
21171 => "000000000000000000000000",
21172 => "000000000000000000000000",
21173 => "000000000000000000000000",
21174 => "000000000000000000000000",
21175 => "000000000000000000000000",
21176 => "000000000000000000000000",
21177 => "000000000000000000000000",
21178 => "000000000000000000000000",
21179 => "000000000000000000000000",
21180 => "001001000010010000100100",
21181 => "010000110100001101000011",
21182 => "010000110100001101000011",
21183 => "010000110100001101000011",
21184 => "010000110100001101000011",
21185 => "010000110100001101000011",
21186 => "010000110100001101000011",
21187 => "010000110100001101000011",
21188 => "010000110100001101000011",
21189 => "010000110100001101000011",
21190 => "010000110100001101000011",
21191 => "010000110100001101000011",
21192 => "010000110100001101000011",
21193 => "010000110100001101000011",
21194 => "010000110100001101000011",
21195 => "010000110100001101000011",
21196 => "010000110100001101000011",
21197 => "010000110100001101000011",
21198 => "010000110100001101000011",
21199 => "000010110000101100001011",
21200 => "000000000000000000000000",
21201 => "000000000000000000000000",
21202 => "000000000000000000000000",
21203 => "000000000000000000000000",
21204 => "000000000000000000000000",
21205 => "000000000000000000000000",
21206 => "000000000000000000000000",
21207 => "000000000000000000000000",
21208 => "000000000000000000000000",
21209 => "000000000000000000000000",
21210 => "000011110000101100000111",
21211 => "111101101011001001101011",
21212 => "111101101011001001101011",
21213 => "111101101011001001101011",
21214 => "111101101011001001101011",
21215 => "100110100110111101000011",
21216 => "000000000000000000000000",
21217 => "000000000000000000000000",
21218 => "000000000000000000000000",
21219 => "000000000000000000000000",
21220 => "000000000000000000000000",
21221 => "000000000000000000000000",
21222 => "010101010011110100100101",
21223 => "111101101011001001101011",
21224 => "111101101011001001101011",
21225 => "000000000000000000000000",
21226 => "000000000000000000000000",
21227 => "000000000000000000000000",
21228 => "000000000000000000000000",
21229 => "000000000000000000000000",
21230 => "000000000000000000000000",
21231 => "000000000000000000000000",
21232 => "000000000000000000000000",
21233 => "000000000000000000000000",
21234 => "000000000000000000000000",
21235 => "000000000000000000000000",
21236 => "000000000000000000000000",
21237 => "000000000000000000000000",
21238 => "000000000000000000000000",
21239 => "010000100100001001000010",
21240 => "010000110100001101000011",
21241 => "010000110100001101000011",
21242 => "010000110100001101000011",
21243 => "010000110100001101000011",
21244 => "010000110100001101000011",
21245 => "010000110100001101000011",
21246 => "010000110100001101000011",
21247 => "010000110100001101000011",
21248 => "010000110100001101000011",
21249 => "010000110100001101000011",
21250 => "010000110100001101000011",
21251 => "010000110100001101000011",
21252 => "010000110100001101000011",
21253 => "010000110100001101000011",
21254 => "010000110100001101000011",
21255 => "010000110100001101000011",
21256 => "010000110100001101000011",
21257 => "001101100011011000110110",
21258 => "000000000000000000000000",
21259 => "000000000000000000000000",
21260 => "000000000000000000000000",
21261 => "000000000000000000000000",
21262 => "000000000000000000000000",
21263 => "000000000000000000000000",
21264 => "000000000000000000000000",
21265 => "000000000000000000000000",
21266 => "000000000000000000000000",
21267 => "000000000000000000000000",
21268 => "000000000000000000000000",
21269 => "000000000000000000000000",
21270 => "000000000000000000000000",
21271 => "000000000000000000000000",
21272 => "000000000000000000000000",
21273 => "000000000000000000000000",
21274 => "000000000000000000000000",
21275 => "000000000000000000000000",
21276 => "000000000000000000000000",
21277 => "000000000000000000000000",
21278 => "000000000000000000000000",
21279 => "000000000000000000000000",
21280 => "000000000000000000000000",
21281 => "000000000000000000000000",
21282 => "000000000000000000000000",
21283 => "000000000000000000000000",
21284 => "000000000000000000000000",
21285 => "000000000000000000000000",
21286 => "000000000000000000000000",
21287 => "000000000000000000000000",
21288 => "000000000000000000000000",
21289 => "000000000000000000000000",
21290 => "000000000000000000000000",
21291 => "000000000000000000000000",
21292 => "000000000000000000000000",
21293 => "000000000000000000000000",
21294 => "000000000000000000000000",
21295 => "000000000000000000000000",
21296 => "000000000000000000000000",
21297 => "000000000000000000000000",
21298 => "000000000000000000000000",
21299 => "000000000000000000000000",
21300 => "000000000000000000000000",
21301 => "000000000000000000000000",
21302 => "000000000000000000000000",
21303 => "000000000000000000000000",
21304 => "000000000000000000000000",
21305 => "000000000000000000000000",
21306 => "000000000000000000000000",
21307 => "000000000000000000000000",
21308 => "000000000000000000000000",
21309 => "000000000000000000000000",
21310 => "000000000000000000000000",
21311 => "000000000000000000000000",
21312 => "000000000000000000000000",
21313 => "000000000000000000000000",
21314 => "000000000000000000000000",
21315 => "000000000000000000000000",
21316 => "000000000000000000000000",
21317 => "000000000000000000000000",
21318 => "000000000000000000000000",
21319 => "000000000000000000000000",
21320 => "000000000000000000000000",
21321 => "000000000000000000000000",
21322 => "000000000000000000000000",
21323 => "000000000000000000000000",
21324 => "000000000000000000000000",
21325 => "000000000000000000000000",
21326 => "000000000000000000000000",
21327 => "000000000000000000000000",
21328 => "000000000000000000000000",
21329 => "000000000000000000000000",
21330 => "001000100010001000100010",
21331 => "010000010100000101000001",
21332 => "010000010100000101000001",
21333 => "010000110100001101000011",
21334 => "010000110100001101000011",
21335 => "010000110100001101000011",
21336 => "010000110100001101000011",
21337 => "010000110100001101000011",
21338 => "010000110100001101000011",
21339 => "010000110100001101000011",
21340 => "010000110100001101000011",
21341 => "010000110100001101000011",
21342 => "010000010100000101000001",
21343 => "010000010100000101000001",
21344 => "010000010100000101000001",
21345 => "010000010100000101000001",
21346 => "010000010100000101000001",
21347 => "010000010100000101000001",
21348 => "010000010100000101000001",
21349 => "000010110000101100001011",
21350 => "000000000000000000000000",
21351 => "000000000000000000000000",
21352 => "000000000000000000000000",
21353 => "000000000000000000000000",
21354 => "000000000000000000000000",
21355 => "000000000000000000000000",
21356 => "000000000000000000000000",
21357 => "000000000000000000000000",
21358 => "000000000000000000000000",
21359 => "000000000000000000000000",
21360 => "000011110000101100000110",
21361 => "111011101010110001101000",
21362 => "111011101010110001101000",
21363 => "111101001011000001101010",
21364 => "111101101011001001101011",
21365 => "100110100110111101000011",
21366 => "000000000000000000000000",
21367 => "000000000000000000000000",
21368 => "000000000000000000000000",
21369 => "000000000000000000000000",
21370 => "000000000000000000000000",
21371 => "000000000000000000000000",
21372 => "010101010011110100100101",
21373 => "111101101011001001101011",
21374 => "111101101011001001101011",
21375 => "000010000000011000000011",
21376 => "000010000000011000000011",
21377 => "000000110000001000000001",
21378 => "000000000000000000000000",
21379 => "000000000000000000000000",
21380 => "000000000000000000000000",
21381 => "000000000000000000000000",
21382 => "000000000000000000000000",
21383 => "000000000000000000000000",
21384 => "000000000000000000000000",
21385 => "000000000000000000000000",
21386 => "000000000000000000000000",
21387 => "000000000000000000000000",
21388 => "000000000000000000000000",
21389 => "010000000100000001000000",
21390 => "010000010100000101000001",
21391 => "010000010100000101000001",
21392 => "010000010100000101000001",
21393 => "010000010100000101000001",
21394 => "010000010100000101000001",
21395 => "010000010100000101000001",
21396 => "010000110100001101000011",
21397 => "010000110100001101000011",
21398 => "010000110100001101000011",
21399 => "010000110100001101000011",
21400 => "010000110100001101000011",
21401 => "010000110100001101000011",
21402 => "010000110100001101000011",
21403 => "010000110100001101000011",
21404 => "010000110100001101000011",
21405 => "010000100100001001000010",
21406 => "010000010100000101000001",
21407 => "001101010011010100110101",
21408 => "000000000000000000000000",
21409 => "000000000000000000000000",
21410 => "000000000000000000000000",
21411 => "000000000000000000000000",
21412 => "000000000000000000000000",
21413 => "000000000000000000000000",
21414 => "000000000000000000000000",
21415 => "000000000000000000000000",
21416 => "000000000000000000000000",
21417 => "000000000000000000000000",
21418 => "000000000000000000000000",
21419 => "000000000000000000000000",
21420 => "000000000000000000000000",
21421 => "000000000000000000000000",
21422 => "000000000000000000000000",
21423 => "000000000000000000000000",
21424 => "000000000000000000000000",
21425 => "000000000000000000000000",
21426 => "000000000000000000000000",
21427 => "000000000000000000000000",
21428 => "000000000000000000000000",
21429 => "000000000000000000000000",
21430 => "000000000000000000000000",
21431 => "000000000000000000000000",
21432 => "000000000000000000000000",
21433 => "000000000000000000000000",
21434 => "000000000000000000000000",
21435 => "000000000000000000000000",
21436 => "000000000000000000000000",
21437 => "000000000000000000000000",
21438 => "000000000000000000000000",
21439 => "000000000000000000000000",
21440 => "000000000000000000000000",
21441 => "000000000000000000000000",
21442 => "000000000000000000000000",
21443 => "000000000000000000000000",
21444 => "000000000000000000000000",
21445 => "000000000000000000000000",
21446 => "000000000000000000000000",
21447 => "000000000000000000000000",
21448 => "000000000000000000000000",
21449 => "000000000000000000000000",
21450 => "000000000000000000000000",
21451 => "000000000000000000000000",
21452 => "000000000000000000000000",
21453 => "000000000000000000000000",
21454 => "000000000000000000000000",
21455 => "000000000000000000000000",
21456 => "000000000000000000000000",
21457 => "000000000000000000000000",
21458 => "000000000000000000000000",
21459 => "000000000000000000000000",
21460 => "000000000000000000000000",
21461 => "000000000000000000000000",
21462 => "000000000000000000000000",
21463 => "000000000000000000000000",
21464 => "000000000000000000000000",
21465 => "000000000000000000000000",
21466 => "000000000000000000000000",
21467 => "000000000000000000000000",
21468 => "000000000000000000000000",
21469 => "000000000000000000000000",
21470 => "000000000000000000000000",
21471 => "000000000000000000000000",
21472 => "000000000000000000000000",
21473 => "000000000000000000000000",
21474 => "000000000000000000000000",
21475 => "000000000000000000000000",
21476 => "000000000000000000000000",
21477 => "000000000000000000000000",
21478 => "000000000000000000000000",
21479 => "000000000000000000000000",
21480 => "000000000000000000000000",
21481 => "000000000000000000000000",
21482 => "000011010000110100001101",
21483 => "010000110100001101000011",
21484 => "010000110100001101000011",
21485 => "010000110100001101000011",
21486 => "010000110100001101000011",
21487 => "010000110100001101000011",
21488 => "010000110100001101000011",
21489 => "010000110100001101000011",
21490 => "010000110100001101000011",
21491 => "010000110100001101000011",
21492 => "000010000000100000001000",
21493 => "000000000000000000000000",
21494 => "000000000000000000000000",
21495 => "000000000000000000000000",
21496 => "000000000000000000000000",
21497 => "000000000000000000000000",
21498 => "000000000000000000000000",
21499 => "000000000000000000000000",
21500 => "000000000000000000000000",
21501 => "000000000000000000000000",
21502 => "000000000000000000000000",
21503 => "000000000000000000000000",
21504 => "000000000000000000000000",
21505 => "000000000000000000000000",
21506 => "000000000000000000000000",
21507 => "000000000000000000000000",
21508 => "000000000000000000000000",
21509 => "000000000000000000000000",
21510 => "000000000000000000000000",
21511 => "000000000000000000000000",
21512 => "000000000000000000000000",
21513 => "101101001000001001001110",
21514 => "111101101011001001101011",
21515 => "100110100110111101000011",
21516 => "000000000000000000000000",
21517 => "000000000000000000000000",
21518 => "000000000000000000000000",
21519 => "000000000000000000000000",
21520 => "000000000000000000000000",
21521 => "000000000000000000000000",
21522 => "010101010011110100100101",
21523 => "111101101011001001101011",
21524 => "111101101011001001101011",
21525 => "111101101011001001101011",
21526 => "111101101011001001101011",
21527 => "010101010011110100100101",
21528 => "000000000000000000000000",
21529 => "000000000000000000000000",
21530 => "000000000000000000000000",
21531 => "000000000000000000000000",
21532 => "000000000000000000000000",
21533 => "000000000000000000000000",
21534 => "000000000000000000000000",
21535 => "000000000000000000000000",
21536 => "000000000000000000000000",
21537 => "000000000000000000000000",
21538 => "000000000000000000000000",
21539 => "000000000000000000000000",
21540 => "000000000000000000000000",
21541 => "000000000000000000000000",
21542 => "000000000000000000000000",
21543 => "000000000000000000000000",
21544 => "000000000000000000000000",
21545 => "000000000000000000000000",
21546 => "010000010100000101000001",
21547 => "010000110100001101000011",
21548 => "010000110100001101000011",
21549 => "010000110100001101000011",
21550 => "010000110100001101000011",
21551 => "010000110100001101000011",
21552 => "010000110100001101000011",
21553 => "010000110100001101000011",
21554 => "010000110100001101000011",
21555 => "000111110001111100011111",
21556 => "000000000000000000000000",
21557 => "000000000000000000000000",
21558 => "000000000000000000000000",
21559 => "000000000000000000000000",
21560 => "000000000000000000000000",
21561 => "000000000000000000000000",
21562 => "000000000000000000000000",
21563 => "000000000000000000000000",
21564 => "000000000000000000000000",
21565 => "000000000000000000000000",
21566 => "000000000000000000000000",
21567 => "000000000000000000000000",
21568 => "000000000000000000000000",
21569 => "000000000000000000000000",
21570 => "000000000000000000000000",
21571 => "000000000000000000000000",
21572 => "000000000000000000000000",
21573 => "000000000000000000000000",
21574 => "000000000000000000000000",
21575 => "000000000000000000000000",
21576 => "000000000000000000000000",
21577 => "000000000000000000000000",
21578 => "000000000000000000000000",
21579 => "000000000000000000000000",
21580 => "000000000000000000000000",
21581 => "000000000000000000000000",
21582 => "000000000000000000000000",
21583 => "000000000000000000000000",
21584 => "000000000000000000000000",
21585 => "000000000000000000000000",
21586 => "000000000000000000000000",
21587 => "000000000000000000000000",
21588 => "000000000000000000000000",
21589 => "000000000000000000000000",
21590 => "000000000000000000000000",
21591 => "000000000000000000000000",
21592 => "000000000000000000000000",
21593 => "000000000000000000000000",
21594 => "000000000000000000000000",
21595 => "000000000000000000000000",
21596 => "000000000000000000000000",
21597 => "000000000000000000000000",
21598 => "000000000000000000000000",
21599 => "000000000000000000000000",
21600 => "000000000000000000000000",
21601 => "000000000000000000000000",
21602 => "000000000000000000000000",
21603 => "000000000000000000000000",
21604 => "000000000000000000000000",
21605 => "000000000000000000000000",
21606 => "000000000000000000000000",
21607 => "000000000000000000000000",
21608 => "000000000000000000000000",
21609 => "000000000000000000000000",
21610 => "000000000000000000000000",
21611 => "000000000000000000000000",
21612 => "000000000000000000000000",
21613 => "000000000000000000000000",
21614 => "000000000000000000000000",
21615 => "000000000000000000000000",
21616 => "000000000000000000000000",
21617 => "000000000000000000000000",
21618 => "000000000000000000000000",
21619 => "000000000000000000000000",
21620 => "000000000000000000000000",
21621 => "000000000000000000000000",
21622 => "000000000000000000000000",
21623 => "000000000000000000000000",
21624 => "000000000000000000000000",
21625 => "000000000000000000000000",
21626 => "000000000000000000000000",
21627 => "000000000000000000000000",
21628 => "000000000000000000000000",
21629 => "000000000000000000000000",
21630 => "000000000000000000000000",
21631 => "000000000000000000000000",
21632 => "000011010000110100001101",
21633 => "010000110100001101000011",
21634 => "010000110100001101000011",
21635 => "010000110100001101000011",
21636 => "010000110100001101000011",
21637 => "010000110100001101000011",
21638 => "010000110100001101000011",
21639 => "010000110100001101000011",
21640 => "010000110100001101000011",
21641 => "010000110100001101000011",
21642 => "000010000000100000001000",
21643 => "000000000000000000000000",
21644 => "000000000000000000000000",
21645 => "000000000000000000000000",
21646 => "000000000000000000000000",
21647 => "000000000000000000000000",
21648 => "000000000000000000000000",
21649 => "000000000000000000000000",
21650 => "000000000000000000000000",
21651 => "000000000000000000000000",
21652 => "000000000000000000000000",
21653 => "000000000000000000000000",
21654 => "000000000000000000000000",
21655 => "000000000000000000000000",
21656 => "000000000000000000000000",
21657 => "000000000000000000000000",
21658 => "000000000000000000000000",
21659 => "000000000000000000000000",
21660 => "000000000000000000000000",
21661 => "000000000000000000000000",
21662 => "000000000000000000000000",
21663 => "101101001000001001001110",
21664 => "111101101011001001101011",
21665 => "100110100110111101000011",
21666 => "000000000000000000000000",
21667 => "000000000000000000000000",
21668 => "000000000000000000000000",
21669 => "000000000000000000000000",
21670 => "000000000000000000000000",
21671 => "000000000000000000000000",
21672 => "010101010011110100100101",
21673 => "111101101011001001101011",
21674 => "111101101011001001101011",
21675 => "111101101011001001101011",
21676 => "111101101011001001101011",
21677 => "010101010011110100100101",
21678 => "000000000000000000000000",
21679 => "000000000000000000000000",
21680 => "000000000000000000000000",
21681 => "000000000000000000000000",
21682 => "000000000000000000000000",
21683 => "000000000000000000000000",
21684 => "000000000000000000000000",
21685 => "000000000000000000000000",
21686 => "000000000000000000000000",
21687 => "000000000000000000000000",
21688 => "000000000000000000000000",
21689 => "000000000000000000000000",
21690 => "000000000000000000000000",
21691 => "000000000000000000000000",
21692 => "000000000000000000000000",
21693 => "000000000000000000000000",
21694 => "000000000000000000000000",
21695 => "000000000000000000000000",
21696 => "010000010100000101000001",
21697 => "010000110100001101000011",
21698 => "010000110100001101000011",
21699 => "010000110100001101000011",
21700 => "010000110100001101000011",
21701 => "010000110100001101000011",
21702 => "010000110100001101000011",
21703 => "010000110100001101000011",
21704 => "010000110100001101000011",
21705 => "000111110001111100011111",
21706 => "000000000000000000000000",
21707 => "000000000000000000000000",
21708 => "000000000000000000000000",
21709 => "000000000000000000000000",
21710 => "000000000000000000000000",
21711 => "000000000000000000000000",
21712 => "000000000000000000000000",
21713 => "000000000000000000000000",
21714 => "000000000000000000000000",
21715 => "000000000000000000000000",
21716 => "000000000000000000000000",
21717 => "000000000000000000000000",
21718 => "000000000000000000000000",
21719 => "000000000000000000000000",
21720 => "000000000000000000000000",
21721 => "000000000000000000000000",
21722 => "000000000000000000000000",
21723 => "000000000000000000000000",
21724 => "000000000000000000000000",
21725 => "000000000000000000000000",
21726 => "000000000000000000000000",
21727 => "000000000000000000000000",
21728 => "000000000000000000000000",
21729 => "000000000000000000000000",
21730 => "000000000000000000000000",
21731 => "000000000000000000000000",
21732 => "000000000000000000000000",
21733 => "000000000000000000000000",
21734 => "000000000000000000000000",
21735 => "000000000000000000000000",
21736 => "000000000000000000000000",
21737 => "000000000000000000000000",
21738 => "000000000000000000000000",
21739 => "000000000000000000000000",
21740 => "000000000000000000000000",
21741 => "000000000000000000000000",
21742 => "000000000000000000000000",
21743 => "000000000000000000000000",
21744 => "000000000000000000000000",
21745 => "000000000000000000000000",
21746 => "000000000000000000000000",
21747 => "000000000000000000000000",
21748 => "000000000000000000000000",
21749 => "000000000000000000000000",
21750 => "000000000000000000000000",
21751 => "000000000000000000000000",
21752 => "000000000000000000000000",
21753 => "000000000000000000000000",
21754 => "000000000000000000000000",
21755 => "000000000000000000000000",
21756 => "000000000000000000000000",
21757 => "000000000000000000000000",
21758 => "000000000000000000000000",
21759 => "000000000000000000000000",
21760 => "000000000000000000000000",
21761 => "000000000000000000000000",
21762 => "000000000000000000000000",
21763 => "000000000000000000000000",
21764 => "000000000000000000000000",
21765 => "000000000000000000000000",
21766 => "000000000000000000000000",
21767 => "000000000000000000000000",
21768 => "000000000000000000000000",
21769 => "000000000000000000000000",
21770 => "000000000000000000000000",
21771 => "000000000000000000000000",
21772 => "000000000000000000000000",
21773 => "000000000000000000000000",
21774 => "000000000000000000000000",
21775 => "000000000000000000000000",
21776 => "000000000000000000000000",
21777 => "000000000000000000000000",
21778 => "000000000000000000000000",
21779 => "000000000000000000000000",
21780 => "000000000000000000000000",
21781 => "000000000000000000000000",
21782 => "000011010000110100001101",
21783 => "010000110100001101000011",
21784 => "010000110100001101000011",
21785 => "010000110100001101000011",
21786 => "010000110100001101000011",
21787 => "001011000010110000101100",
21788 => "000101010001010100010101",
21789 => "000101010001010100010101",
21790 => "000101010001010100010101",
21791 => "000101010001010100010101",
21792 => "000000110000001100000011",
21793 => "000000000000000000000000",
21794 => "000000000000000000000000",
21795 => "000000000000000000000000",
21796 => "000000000000000000000000",
21797 => "000000000000000000000000",
21798 => "000000000000000000000000",
21799 => "000000000000000000000000",
21800 => "000000000000000000000000",
21801 => "000000000000000000000000",
21802 => "000000000000000000000000",
21803 => "000000000000000000000000",
21804 => "000000000000000000000000",
21805 => "000000000000000000000000",
21806 => "000000000000000000000000",
21807 => "000000000000000000000000",
21808 => "000000000000000000000000",
21809 => "000000000000000000000000",
21810 => "000010110000100000000101",
21811 => "101010010111101001001010",
21812 => "101010010111101001001010",
21813 => "011001100100101000101100",
21814 => "010011010011100000100001",
21815 => "001100000010001100010101",
21816 => "000000000000000000000000",
21817 => "000000000000000000000000",
21818 => "000000000000000000000000",
21819 => "000000000000000000000000",
21820 => "000000000000000000000000",
21821 => "000000000000000000000000",
21822 => "000110100001001100001011",
21823 => "010011010011100000100001",
21824 => "010011010011100000100001",
21825 => "111101101011001001101011",
21826 => "111101101011001001101011",
21827 => "010101010011110100100101",
21828 => "000000000000000000000000",
21829 => "000000000000000000000000",
21830 => "000000000000000000000000",
21831 => "000000000000000000000000",
21832 => "000000000000000000000000",
21833 => "000000000000000000000000",
21834 => "000000000000000000000000",
21835 => "000000000000000000000000",
21836 => "000000000000000000000000",
21837 => "000000000000000000000000",
21838 => "000000000000000000000000",
21839 => "000000000000000000000000",
21840 => "000000000000000000000000",
21841 => "000000000000000000000000",
21842 => "000000000000000000000000",
21843 => "000000000000000000000000",
21844 => "000000000000000000000000",
21845 => "000000000000000000000000",
21846 => "000101000001010000010100",
21847 => "000101010001010100010101",
21848 => "000101010001010100010101",
21849 => "000101010001010100010101",
21850 => "000111110001111100011111",
21851 => "010000110100001101000011",
21852 => "010000110100001101000011",
21853 => "010000110100001101000011",
21854 => "010000110100001101000011",
21855 => "000111110001111100011111",
21856 => "000000000000000000000000",
21857 => "000000000000000000000000",
21858 => "000000000000000000000000",
21859 => "000000000000000000000000",
21860 => "000000000000000000000000",
21861 => "000000000000000000000000",
21862 => "000000000000000000000000",
21863 => "000000000000000000000000",
21864 => "000000000000000000000000",
21865 => "000000000000000000000000",
21866 => "000000000000000000000000",
21867 => "000000000000000000000000",
21868 => "000000000000000000000000",
21869 => "000000000000000000000000",
21870 => "000000000000000000000000",
21871 => "000000000000000000000000",
21872 => "000000000000000000000000",
21873 => "000000000000000000000000",
21874 => "000000000000000000000000",
21875 => "000000000000000000000000",
21876 => "000000000000000000000000",
21877 => "000000000000000000000000",
21878 => "000000000000000000000000",
21879 => "000000000000000000000000",
21880 => "000000000000000000000000",
21881 => "000000000000000000000000",
21882 => "000000000000000000000000",
21883 => "000000000000000000000000",
21884 => "000000000000000000000000",
21885 => "000000000000000000000000",
21886 => "000000000000000000000000",
21887 => "000000000000000000000000",
21888 => "000000000000000000000000",
21889 => "000000000000000000000000",
21890 => "000000000000000000000000",
21891 => "000000000000000000000000",
21892 => "000000000000000000000000",
21893 => "000000000000000000000000",
21894 => "000000000000000000000000",
21895 => "000000000000000000000000",
21896 => "000000000000000000000000",
21897 => "000000000000000000000000",
21898 => "000000000000000000000000",
21899 => "000000000000000000000000",
21900 => "000000000000000000000000",
21901 => "000000000000000000000000",
21902 => "000000000000000000000000",
21903 => "000000000000000000000000",
21904 => "000000000000000000000000",
21905 => "000000000000000000000000",
21906 => "000000000000000000000000",
21907 => "000000000000000000000000",
21908 => "000000000000000000000000",
21909 => "000000000000000000000000",
21910 => "000000000000000000000000",
21911 => "000000000000000000000000",
21912 => "000000000000000000000000",
21913 => "000000000000000000000000",
21914 => "000000000000000000000000",
21915 => "000000000000000000000000",
21916 => "000000000000000000000000",
21917 => "000000000000000000000000",
21918 => "000000000000000000000000",
21919 => "000000000000000000000000",
21920 => "000000000000000000000000",
21921 => "000000000000000000000000",
21922 => "000000000000000000000000",
21923 => "000000000000000000000000",
21924 => "000000000000000000000000",
21925 => "000000000000000000000000",
21926 => "000000000000000000000000",
21927 => "000000000000000000000000",
21928 => "000000000000000000000000",
21929 => "000000000000000000000000",
21930 => "000000000000000000000000",
21931 => "000000000000000000000000",
21932 => "000011010000110100001101",
21933 => "010000110100001101000011",
21934 => "010000110100001101000011",
21935 => "010000110100001101000011",
21936 => "010000110100001101000011",
21937 => "001000100010001000100010",
21938 => "000000000000000000000000",
21939 => "000000000000000000000000",
21940 => "000000000000000000000000",
21941 => "000000000000000000000000",
21942 => "000000000000000000000000",
21943 => "000000000000000000000000",
21944 => "000000000000000000000000",
21945 => "000000000000000000000000",
21946 => "000000000000000000000000",
21947 => "000000000000000000000000",
21948 => "000000000000000000000000",
21949 => "000000000000000000000000",
21950 => "000000000000000000000000",
21951 => "000000000000000000000000",
21952 => "000000000000000000000000",
21953 => "000000000000000000000000",
21954 => "000000000000000000000000",
21955 => "000000000000000000000000",
21956 => "000000000000000000000000",
21957 => "000000000000000000000000",
21958 => "000000000000000000000000",
21959 => "000000000000000000000000",
21960 => "000011110000101100000111",
21961 => "111101101011001001101011",
21962 => "111101101011001001101011",
21963 => "010000100011000000011101",
21964 => "000000000000000000000000",
21965 => "000000000000000000000000",
21966 => "000000000000000000000000",
21967 => "000000000000000000000000",
21968 => "000000000000000000000000",
21969 => "000000000000000000000000",
21970 => "000000000000000000000000",
21971 => "000000000000000000000000",
21972 => "000000000000000000000000",
21973 => "000000000000000000000000",
21974 => "000000000000000000000000",
21975 => "111101101011001001101011",
21976 => "111101101011001001101011",
21977 => "010101010011110100100101",
21978 => "000000000000000000000000",
21979 => "000000000000000000000000",
21980 => "000000000000000000000000",
21981 => "000000000000000000000000",
21982 => "000000000000000000000000",
21983 => "000000000000000000000000",
21984 => "000000000000000000000000",
21985 => "000000000000000000000000",
21986 => "000000000000000000000000",
21987 => "000000000000000000000000",
21988 => "000000000000000000000000",
21989 => "000000000000000000000000",
21990 => "000000000000000000000000",
21991 => "000000000000000000000000",
21992 => "000000000000000000000000",
21993 => "000000000000000000000000",
21994 => "000000000000000000000000",
21995 => "000000000000000000000000",
21996 => "000000000000000000000000",
21997 => "000000000000000000000000",
21998 => "000000000000000000000000",
21999 => "000000000000000000000000",
22000 => "000011110000111100001111",
22001 => "010000110100001101000011",
22002 => "010000110100001101000011",
22003 => "010000110100001101000011",
22004 => "010000110100001101000011",
22005 => "000111110001111100011111",
22006 => "000000000000000000000000",
22007 => "000000000000000000000000",
22008 => "000000000000000000000000",
22009 => "000000000000000000000000",
22010 => "000000000000000000000000",
22011 => "000000000000000000000000",
22012 => "000000000000000000000000",
22013 => "000000000000000000000000",
22014 => "000000000000000000000000",
22015 => "000000000000000000000000",
22016 => "000000000000000000000000",
22017 => "000000000000000000000000",
22018 => "000000000000000000000000",
22019 => "000000000000000000000000",
22020 => "000000000000000000000000",
22021 => "000000000000000000000000",
22022 => "000000000000000000000000",
22023 => "000000000000000000000000",
22024 => "000000000000000000000000",
22025 => "000000000000000000000000",
22026 => "000000000000000000000000",
22027 => "000000000000000000000000",
22028 => "000000000000000000000000",
22029 => "000000000000000000000000",
22030 => "000000000000000000000000",
22031 => "000000000000000000000000",
22032 => "000000000000000000000000",
22033 => "000000000000000000000000",
22034 => "000000000000000000000000",
22035 => "000000000000000000000000",
22036 => "000000000000000000000000",
22037 => "000000000000000000000000",
22038 => "000000000000000000000000",
22039 => "000000000000000000000000",
22040 => "000000000000000000000000",
22041 => "000000000000000000000000",
22042 => "000000000000000000000000",
22043 => "000000000000000000000000",
22044 => "000000000000000000000000",
22045 => "000000000000000000000000",
22046 => "000000000000000000000000",
22047 => "000000000000000000000000",
22048 => "000000000000000000000000",
22049 => "000000000000000000000000",
22050 => "000000000000000000000000",
22051 => "000000000000000000000000",
22052 => "000000000000000000000000",
22053 => "000000000000000000000000",
22054 => "000000000000000000000000",
22055 => "000000000000000000000000",
22056 => "000000000000000000000000",
22057 => "000000000000000000000000",
22058 => "000000000000000000000000",
22059 => "000000000000000000000000",
22060 => "000000000000000000000000",
22061 => "000000000000000000000000",
22062 => "000000000000000000000000",
22063 => "000000000000000000000000",
22064 => "000000000000000000000000",
22065 => "000000000000000000000000",
22066 => "000000000000000000000000",
22067 => "000000000000000000000000",
22068 => "000000000000000000000000",
22069 => "000000000000000000000000",
22070 => "000000000000000000000000",
22071 => "000000000000000000000000",
22072 => "000000000000000000000000",
22073 => "000000000000000000000000",
22074 => "000000000000000000000000",
22075 => "000000000000000000000000",
22076 => "000000000000000000000000",
22077 => "000000000000000000000000",
22078 => "000000000000000000000000",
22079 => "000000000000000000000000",
22080 => "000000000000000000000000",
22081 => "000000000000000000000000",
22082 => "000010000000100000001000",
22083 => "001011000010110000101100",
22084 => "001011000010110000101100",
22085 => "001011000010110000101100",
22086 => "001011000010110000101100",
22087 => "000101100001011000010110",
22088 => "000000000000000000000000",
22089 => "000000000000000000000000",
22090 => "000000000000000000000000",
22091 => "000000000000000000000000",
22092 => "000000000000000000000000",
22093 => "000000000000000000000000",
22094 => "000000000000000000000000",
22095 => "000000000000000000000000",
22096 => "000000000000000000000000",
22097 => "000000000000000000000000",
22098 => "000000000000000000000000",
22099 => "000000000000000000000000",
22100 => "000000000000000000000000",
22101 => "000000000000000000000000",
22102 => "000000000000000000000000",
22103 => "000000000000000000000000",
22104 => "000000000000000000000000",
22105 => "000000000000000000000000",
22106 => "000000000000000000000000",
22107 => "000000000000000000000000",
22108 => "000000000000000000000000",
22109 => "000000000000000000000000",
22110 => "000010100000011100000100",
22111 => "101000010111010101000110",
22112 => "101000010111010101000110",
22113 => "001011000010000000010011",
22114 => "000000000000000000000000",
22115 => "000000000000000000000000",
22116 => "000000000000000000000000",
22117 => "000000000000000000000000",
22118 => "000000000000000000000000",
22119 => "000000000000000000000000",
22120 => "000000000000000000000000",
22121 => "000000000000000000000000",
22122 => "000000000000000000000000",
22123 => "000000000000000000000000",
22124 => "000000000000000000000000",
22125 => "101000010111010101000110",
22126 => "101000010111010101000110",
22127 => "001101110010100000011000",
22128 => "000000000000000000000000",
22129 => "000000000000000000000000",
22130 => "000000000000000000000000",
22131 => "000000000000000000000000",
22132 => "000000000000000000000000",
22133 => "000000000000000000000000",
22134 => "000000000000000000000000",
22135 => "000000000000000000000000",
22136 => "000000000000000000000000",
22137 => "000000000000000000000000",
22138 => "000000000000000000000000",
22139 => "000000000000000000000000",
22140 => "000000000000000000000000",
22141 => "000000000000000000000000",
22142 => "000000000000000000000000",
22143 => "000000000000000000000000",
22144 => "000000000000000000000000",
22145 => "000000000000000000000000",
22146 => "000000000000000000000000",
22147 => "000000000000000000000000",
22148 => "000000000000000000000000",
22149 => "000000000000000000000000",
22150 => "000010100000101000001010",
22151 => "001011000010110000101100",
22152 => "001011000010110000101100",
22153 => "001011000010110000101100",
22154 => "001011000010110000101100",
22155 => "000101010001010100010101",
22156 => "000000000000000000000000",
22157 => "000000000000000000000000",
22158 => "000000000000000000000000",
22159 => "000000000000000000000000",
22160 => "000000000000000000000000",
22161 => "000000000000000000000000",
22162 => "000000000000000000000000",
22163 => "000000000000000000000000",
22164 => "000000000000000000000000",
22165 => "000000000000000000000000",
22166 => "000000000000000000000000",
22167 => "000000000000000000000000",
22168 => "000000000000000000000000",
22169 => "000000000000000000000000",
22170 => "000000000000000000000000",
22171 => "000000000000000000000000",
22172 => "000000000000000000000000",
22173 => "000000000000000000000000",
22174 => "000000000000000000000000",
22175 => "000000000000000000000000",
22176 => "000000000000000000000000",
22177 => "000000000000000000000000",
22178 => "000000000000000000000000",
22179 => "000000000000000000000000",
22180 => "000000000000000000000000",
22181 => "000000000000000000000000",
22182 => "000000000000000000000000",
22183 => "000000000000000000000000",
22184 => "000000000000000000000000",
22185 => "000000000000000000000000",
22186 => "000000000000000000000000",
22187 => "000000000000000000000000",
22188 => "000000000000000000000000",
22189 => "000000000000000000000000",
22190 => "000000000000000000000000",
22191 => "000000000000000000000000",
22192 => "000000000000000000000000",
22193 => "000000000000000000000000",
22194 => "000000000000000000000000",
22195 => "000000000000000000000000",
22196 => "000000000000000000000000",
22197 => "000000000000000000000000",
22198 => "000000000000000000000000",
22199 => "000000000000000000000000",
22200 => "000000000000000000000000",
22201 => "000000000000000000000000",
22202 => "000000000000000000000000",
22203 => "000000000000000000000000",
22204 => "000000000000000000000000",
22205 => "000000000000000000000000",
22206 => "000000000000000000000000",
22207 => "000000000000000000000000",
22208 => "000000000000000000000000",
22209 => "000000000000000000000000",
22210 => "000000000000000000000000",
22211 => "000000000000000000000000",
22212 => "000000000000000000000000",
22213 => "000000000000000000000000",
22214 => "000000000000000000000000",
22215 => "000000000000000000000000",
22216 => "000000000000000000000000",
22217 => "000000000000000000000000",
22218 => "000000000000000000000000",
22219 => "000000000000000000000000",
22220 => "000000000000000000000000",
22221 => "000000000000000000000000",
22222 => "000000000000000000000000",
22223 => "000000000000000000000000",
22224 => "000000000000000000000000",
22225 => "000000000000000000000000",
22226 => "000000000000000000000000",
22227 => "000000000000000000000000",
22228 => "000000000000000000000000",
22229 => "000000000000000000000000",
22230 => "000000000000000000000000",
22231 => "000000000000000000000000",
22232 => "000000000000000000000000",
22233 => "000000000000000000000000",
22234 => "000000000000000000000000",
22235 => "000000000000000000000000",
22236 => "000000000000000000000000",
22237 => "000000000000000000000000",
22238 => "000000000000000000000000",
22239 => "000000000000000000000000",
22240 => "000000000000000000000000",
22241 => "000000000000000000000000",
22242 => "000000000000000000000000",
22243 => "000000000000000000000000",
22244 => "000000000000000000000000",
22245 => "000000000000000000000000",
22246 => "000000000000000000000000",
22247 => "000000000000000000000000",
22248 => "000000000000000000000000",
22249 => "000000000000000000000000",
22250 => "000000000000000000000000",
22251 => "000000000000000000000000",
22252 => "000000000000000000000000",
22253 => "000000000000000000000000",
22254 => "000000000000000000000000",
22255 => "000000000000000000000000",
22256 => "000000000000000000000000",
22257 => "000000000000000000000000",
22258 => "000000000000000000000000",
22259 => "000000000000000000000000",
22260 => "000000000000000000000000",
22261 => "000000000000000000000000",
22262 => "000000000000000000000000",
22263 => "000000000000000000000000",
22264 => "000000000000000000000000",
22265 => "000000000000000000000000",
22266 => "000000000000000000000000",
22267 => "000000000000000000000000",
22268 => "000000000000000000000000",
22269 => "000000000000000000000000",
22270 => "000000000000000000000000",
22271 => "000000000000000000000000",
22272 => "000000000000000000000000",
22273 => "000000000000000000000000",
22274 => "000000000000000000000000",
22275 => "000000000000000000000000",
22276 => "000000000000000000000000",
22277 => "000000000000000000000000",
22278 => "000000000000000000000000",
22279 => "000000000000000000000000",
22280 => "000000000000000000000000",
22281 => "000000000000000000000000",
22282 => "000000000000000000000000",
22283 => "000000000000000000000000",
22284 => "000000000000000000000000",
22285 => "000000000000000000000000",
22286 => "000000000000000000000000",
22287 => "000000000000000000000000",
22288 => "000000000000000000000000",
22289 => "000000000000000000000000",
22290 => "000000000000000000000000",
22291 => "000000000000000000000000",
22292 => "000000000000000000000000",
22293 => "000000000000000000000000",
22294 => "000000000000000000000000",
22295 => "000000000000000000000000",
22296 => "000000000000000000000000",
22297 => "000000000000000000000000",
22298 => "000000000000000000000000",
22299 => "000000000000000000000000",
22300 => "000000000000000000000000",
22301 => "000000000000000000000000",
22302 => "000000000000000000000000",
22303 => "000000000000000000000000",
22304 => "000000000000000000000000",
22305 => "000000000000000000000000",
22306 => "000000000000000000000000",
22307 => "000000000000000000000000",
22308 => "000000000000000000000000",
22309 => "000000000000000000000000",
22310 => "000000000000000000000000",
22311 => "000000000000000000000000",
22312 => "000000000000000000000000",
22313 => "000000000000000000000000",
22314 => "000000000000000000000000",
22315 => "000000000000000000000000",
22316 => "000000000000000000000000",
22317 => "000000000000000000000000",
22318 => "000000000000000000000000",
22319 => "000000000000000000000000",
22320 => "000000000000000000000000",
22321 => "000000000000000000000000",
22322 => "000000000000000000000000",
22323 => "000000000000000000000000",
22324 => "000000000000000000000000",
22325 => "000000000000000000000000",
22326 => "000000000000000000000000",
22327 => "000000000000000000000000",
22328 => "000000000000000000000000",
22329 => "000000000000000000000000",
22330 => "000000000000000000000000",
22331 => "000000000000000000000000",
22332 => "000000000000000000000000",
22333 => "000000000000000000000000",
22334 => "000000000000000000000000",
22335 => "000000000000000000000000",
22336 => "000000000000000000000000",
22337 => "000000000000000000000000",
22338 => "000000000000000000000000",
22339 => "000000000000000000000000",
22340 => "000000000000000000000000",
22341 => "000000000000000000000000",
22342 => "000000000000000000000000",
22343 => "000000000000000000000000",
22344 => "000000000000000000000000",
22345 => "000000000000000000000000",
22346 => "000000000000000000000000",
22347 => "000000000000000000000000",
22348 => "000000000000000000000000",
22349 => "000000000000000000000000",
22350 => "000000000000000000000000",
22351 => "000000000000000000000000",
22352 => "000000000000000000000000",
22353 => "000000000000000000000000",
22354 => "000000000000000000000000",
22355 => "000000000000000000000000",
22356 => "000000000000000000000000",
22357 => "000000000000000000000000",
22358 => "000000000000000000000000",
22359 => "000000000000000000000000",
22360 => "000000000000000000000000",
22361 => "000000000000000000000000",
22362 => "000000000000000000000000",
22363 => "000000000000000000000000",
22364 => "000000000000000000000000",
22365 => "000000000000000000000000",
22366 => "000000000000000000000000",
22367 => "000000000000000000000000",
22368 => "000000000000000000000000",
22369 => "000000000000000000000000",
22370 => "000000000000000000000000",
22371 => "000000000000000000000000",
22372 => "000000000000000000000000",
22373 => "000000000000000000000000",
22374 => "000000000000000000000000",
22375 => "000000000000000000000000",
22376 => "000000000000000000000000",
22377 => "000000000000000000000000",
22378 => "000000000000000000000000",
22379 => "000000000000000000000000",
22380 => "000000000000000000000000",
22381 => "000000000000000000000000",
22382 => "000000000000000000000000",
22383 => "000000000000000000000000",
22384 => "000000000000000000000000",
22385 => "000000000000000000000000",
22386 => "000000000000000000000000",
22387 => "000000000000000000000000",
22388 => "000000000000000000000000",
22389 => "000000000000000000000000",
22390 => "000000000000000000000000",
22391 => "000000000000000000000000",
22392 => "000000000000000000000000",
22393 => "000000000000000000000000",
22394 => "000000000000000000000000",
22395 => "000000000000000000000000",
22396 => "000000000000000000000000",
22397 => "000000000000000000000000",
22398 => "000000000000000000000000",
22399 => "000000000000000000000000",
22400 => "000000000000000000000000",
22401 => "000000000000000000000000",
22402 => "000000000000000000000000",
22403 => "000000000000000000000000",
22404 => "000000000000000000000000",
22405 => "000000000000000000000000",
22406 => "000000000000000000000000",
22407 => "000000000000000000000000",
22408 => "000000000000000000000000",
22409 => "000000000000000000000000",
22410 => "000000000000000000000000",
22411 => "000000000000000000000000",
22412 => "000000000000000000000000",
22413 => "000000000000000000000000",
22414 => "000000000000000000000000",
22415 => "000000000000000000000000",
22416 => "000000000000000000000000",
22417 => "000000000000000000000000",
22418 => "000000000000000000000000",
22419 => "000000000000000000000000",
22420 => "000000000000000000000000",
22421 => "000000000000000000000000",
22422 => "000000000000000000000000",
22423 => "000000000000000000000000",
22424 => "000000000000000000000000",
22425 => "000000000000000000000000",
22426 => "000000000000000000000000",
22427 => "000000000000000000000000",
22428 => "000000000000000000000000",
22429 => "000000000000000000000000",
22430 => "000000000000000000000000",
22431 => "000000000000000000000000",
22432 => "000000000000000000000000",
22433 => "000000000000000000000000",
22434 => "000000000000000000000000",
22435 => "000000000000000000000000",
22436 => "000000000000000000000000",
22437 => "000000000000000000000000",
22438 => "000000000000000000000000",
22439 => "000000000000000000000000",
22440 => "000000000000000000000000",
22441 => "000000000000000000000000",
22442 => "000000000000000000000000",
22443 => "000000000000000000000000",
22444 => "000000000000000000000000",
22445 => "000000000000000000000000",
22446 => "000000000000000000000000",
22447 => "000000000000000000000000",
22448 => "000000000000000000000000",
22449 => "000000000000000000000000",
22450 => "000000000000000000000000",
22451 => "000000000000000000000000",
22452 => "000000000000000000000000",
22453 => "000000000000000000000000",
22454 => "000000000000000000000000",
22455 => "000000000000000000000000",
22456 => "000000000000000000000000",
22457 => "000000000000000000000000",
22458 => "000000000000000000000000",
22459 => "000000000000000000000000",
22460 => "000000000000000000000000",
22461 => "000000000000000000000000",
22462 => "000000000000000000000000",
22463 => "000000000000000000000000",
22464 => "000000000000000000000000",
22465 => "000000000000000000000000",
22466 => "000000000000000000000000",
22467 => "000000000000000000000000",
22468 => "000000000000000000000000",
22469 => "000000000000000000000000",
22470 => "000000000000000000000000",
22471 => "000000000000000000000000",
22472 => "000000000000000000000000",
22473 => "000000000000000000000000",
22474 => "000000000000000000000000",
22475 => "000000000000000000000000",
22476 => "000000000000000000000000",
22477 => "000000000000000000000000",
22478 => "000000000000000000000000",
22479 => "000000000000000000000000",
22480 => "000000000000000000000000",
22481 => "000000000000000000000000",
22482 => "000000000000000000000000",
22483 => "000000000000000000000000",
22484 => "000000000000000000000000",
22485 => "000000000000000000000000",
22486 => "000000000000000000000000",
22487 => "000000000000000000000000",
22488 => "000000000000000000000000",
22489 => "000000000000000000000000",
22490 => "000000000000000000000000",
22491 => "000000000000000000000000",
22492 => "000000000000000000000000",
22493 => "000000000000000000000000",
22494 => "000000000000000000000000",
22495 => "000000000000000000000000",
22496 => "000000000000000000000000",
22497 => "000000000000000000000000",
22498 => "000000000000000000000000",
22499 => "000000000000000000000000"


    );
begin
    data_out <= ROM_Data(to_integer(unsigned(address)));
end architecture Behavioral;