library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;
use ieee.numeric_std.all;

entity creditsComp is
    Port (
        address : in STD_LOGIC_VECTOR(12 downto 0);
        data_out : out STD_LOGIC_VECTOR(23 downto 0)
    );
end entity creditsComp;

architecture Behavioral of creditsComp is
    type ROM_Type is array (0 to 4199) of STD_LOGIC_VECTOR(23 downto 0);
    constant ROM_Data : ROM_Type := (
0 => "000001000000010000000100",
1 => "000001100000011000000110",
2 => "000001100000011000000110",
3 => "000001100000011000000110",
4 => "000001100000011000000110",
5 => "000000100000001000000010",
6 => "000000000000000000000000",
7 => "000000000000000000000000",
8 => "000000000000000000000000",
9 => "000000000000000000000000",
10 => "000000000000000000000000",
11 => "000000000000000000000000",
12 => "000000000000000000000000",
13 => "000000000000000000000000",
14 => "000000000000000000000000",
15 => "000000000000000000000000",
16 => "000000000000000000000000",
17 => "000000000000000000000000",
18 => "000000000000000000000000",
19 => "000000000000000000000000",
20 => "000000000000000000000000",
21 => "000000000000000000000000",
22 => "000000000000000000000000",
23 => "000000000000000000000000",
24 => "000000000000000000000000",
25 => "000000000000000000000000",
26 => "000000000000000000000000",
27 => "000000000000000000000000",
28 => "000000000000000000000000",
29 => "000000000000000000000000",
30 => "000000000000000000000000",
31 => "000000000000000000000000",
32 => "000000110000001100000011",
33 => "000001100000011000000110",
34 => "000001010000010100000101",
35 => "000000100000001000000010",
36 => "000001100000011000000110",
37 => "011010000110100001101000",
38 => "011001110110011101100111",
39 => "000001010000010100000101",
40 => "000000000000000000000000",
41 => "000000000000000000000000",
42 => "000000000000000000000000",
43 => "000000000000000000000000",
44 => "000000000000000000000000",
45 => "000000000000000000000000",
46 => "000000000000000000000000",
47 => "000000000000000000000000",
48 => "000000000000000000000000",
49 => "000000000000000000000000",
50 => "010010110100101101001011",
51 => "011110010111100101111001",
52 => "000100100001001000010010",
53 => "000000000000000000000000",
54 => "000000000000000000000000",
55 => "000000000000000000000000",
56 => "000000000000000000000000",
57 => "000000000000000000000000",
58 => "000000000000000000000000",
59 => "000000000000000000000000",
60 => "000000000000000000000000",
61 => "000000000000000000000000",
62 => "000000000000000000000000",
63 => "000000000000000000000000",
64 => "000000000000000000000000",
65 => "000000000000000000000000",
66 => "000000000000000000000000",
67 => "000000000000000000000000",
68 => "000000000000000000000000",
69 => "000000000000000000000000",
70 => "000000000000000000000000",
71 => "000000000000000000000000",
72 => "000000000000000000000000",
73 => "000000000000000000000000",
74 => "000000000000000000000000",
75 => "000000000000000000000000",
76 => "000000000000000000000000",
77 => "000000000000000000000000",
78 => "000000000000000000000000",
79 => "000000000000000000000000",
80 => "000000000000000000000000",
81 => "000000000000000000000000",
82 => "000000000000000000000000",
83 => "000000000000000000000000",
84 => "000000000000000000000000",
85 => "000000000000000000000000",
86 => "000000000000000000000000",
87 => "000000000000000000000000",
88 => "000000000000000000000000",
89 => "000000000000000000000000",
90 => "000000000000000000000000",
91 => "000000000000000000000000",
92 => "000000000000000000000000",
93 => "000000000000000000000000",
94 => "000000000000000000000000",
95 => "000000000000000000000000",
96 => "000000000000000000000000",
97 => "000000000000000000000000",
98 => "000000000000000000000000",
99 => "000000000000000000000000",
100 => "100110111001101110011011",
101 => "111111111111111111111111",
102 => "111111101111111011111110",
103 => "111110011111100111111001",
104 => "111111111111111111111111",
105 => "011000000110000001100000",
106 => "000000000000000000000000",
107 => "000000000000000000000000",
108 => "000000000000000000000000",
109 => "000000000000000000000000",
110 => "000000000000000000000000",
111 => "000000000000000000000000",
112 => "000000000000000000000000",
113 => "000000000000000000000000",
114 => "000000000000000000000000",
115 => "000000000000000000000000",
116 => "000000000000000000000000",
117 => "000000000000000000000000",
118 => "000000000000000000000000",
119 => "000000000000000000000000",
120 => "000000000000000000000000",
121 => "000000000000000000000000",
122 => "000000000000000000000000",
123 => "000000000000000000000000",
124 => "000000000000000000000000",
125 => "000000000000000000000000",
126 => "000000000000000000000000",
127 => "000000000000000000000000",
128 => "000000000000000000000000",
129 => "000000000000000000000000",
130 => "000000010000000100000001",
131 => "010101100101011001010110",
132 => "110011111100111111001111",
133 => "111101111111011111110111",
134 => "111011111110111111101111",
135 => "101100011011000110110001",
136 => "000111100001111000011110",
137 => "110111101101111011011110",
138 => "110011011100110111001101",
139 => "000100000001000000010000",
140 => "000000000000000000000000",
141 => "000000000000000000000000",
142 => "000000000000000000000000",
143 => "000000000000000000000000",
144 => "000000000000000000000000",
145 => "000000000000000000000000",
146 => "000000000000000000000000",
147 => "000000010000000100000001",
148 => "000000000000000000000000",
149 => "000000000000000000000000",
150 => "101100111011001110110011",
151 => "111010001110100011101000",
152 => "001100000011000000110000",
153 => "000000000000000000000000",
154 => "000000000000000000000000",
155 => "000000000000000000000000",
156 => "000000000000000000000000",
157 => "000000000000000000000000",
158 => "000000000000000000000000",
159 => "000000000000000000000000",
160 => "000000000000000000000000",
161 => "000000000000000000000000",
162 => "000000000000000000000000",
163 => "000000000000000000000000",
164 => "000000000000000000000000",
165 => "000000000000000000000000",
166 => "000000000000000000000000",
167 => "000000000000000000000000",
168 => "000000000000000000000000",
169 => "000000000000000000000000",
170 => "000000000000000000000000",
171 => "000000000000000000000000",
172 => "000000000000000000000000",
173 => "000000000000000000000000",
174 => "000000000000000000000000",
175 => "000000000000000000000000",
176 => "000000000000000000000000",
177 => "000000000000000000000000",
178 => "000000000000000000000000",
179 => "000000000000000000000000",
180 => "000000000000000000000000",
181 => "000000000000000000000000",
182 => "000000000000000000000000",
183 => "000000000000000000000000",
184 => "000000000000000000000000",
185 => "000000000000000000000000",
186 => "000000000000000000000000",
187 => "000000000000000000000000",
188 => "000000000000000000000000",
189 => "000000000000000000000000",
190 => "000000000000000000000000",
191 => "000000000000000000000000",
192 => "000000000000000000000000",
193 => "000000000000000000000000",
194 => "000000000000000000000000",
195 => "000000000000000000000000",
196 => "000000000000000000000000",
197 => "000000000000000000000000",
198 => "000000000000000000000000",
199 => "000000000000000000000000",
200 => "000101110001011100010111",
201 => "111111111111111111111111",
202 => "110011101100111011001110",
203 => "001110110011101100111011",
204 => "110101011101010111010101",
205 => "010110110101101101011011",
206 => "001111010011110100111101",
207 => "100101011001010110010101",
208 => "011100010111000101110001",
209 => "000011000000110000001100",
210 => "010001110100011101000111",
211 => "100110011001100110011001",
212 => "100110011001100110011001",
213 => "010010010100100101001001",
214 => "100110001001100010011000",
215 => "100110011001100110011001",
216 => "001101100011011000110110",
217 => "100110011001100110011001",
218 => "100110011001100110011001",
219 => "100110011001100110011001",
220 => "100101001001010010010100",
221 => "000111010001110100011101",
222 => "001100110011001100110011",
223 => "100000001000000010000000",
224 => "100110011001100110011001",
225 => "011010000110100001101000",
226 => "000010000000100000001000",
227 => "000000000000000000000000",
228 => "000000000000000000000000",
229 => "000000000000000000000000",
230 => "001110010011100100111001",
231 => "111110101111101011111010",
232 => "101010111010101110101011",
233 => "001001000010010000100100",
234 => "101010111010101110101011",
235 => "111100001111000011110000",
236 => "000110010001100100011001",
237 => "001001000010010000100100",
238 => "001011100010111000101110",
239 => "000110110001101100011011",
240 => "100100101001001010010010",
241 => "100110011001100110011001",
242 => "011011100110111001101110",
243 => "100011001000110010001100",
244 => "100110011001100110011001",
245 => "011100000111000001110000",
246 => "100110001001100010011000",
247 => "100011011000110110001101",
248 => "010101010101010101010101",
249 => "011100010111000101110001",
250 => "000110110001101100011011",
251 => "001100010011000100110001",
252 => "000011100000111000001110",
253 => "000000000000000000000000",
254 => "000000000000000000000000",
255 => "000000000000000000000000",
256 => "000000000000000000000000",
257 => "000000000000000000000000",
258 => "000000000000000000000000",
259 => "000000000000000000000000",
260 => "000000000000000000000000",
261 => "000000000000000000000000",
262 => "000000000000000000000000",
263 => "000000000000000000000000",
264 => "000000000000000000000000",
265 => "000000000000000000000000",
266 => "000000000000000000000000",
267 => "000000000000000000000000",
268 => "000000000000000000000000",
269 => "000000000000000000000000",
270 => "000000000000000000000000",
271 => "000000000000000000000000",
272 => "000000000000000000000000",
273 => "000000000000000000000000",
274 => "000000000000000000000000",
275 => "000000000000000000000000",
276 => "000000000000000000000000",
277 => "000000000000000000000000",
278 => "000000000000000000000000",
279 => "000000000000000000000000",
280 => "000000000000000000000000",
281 => "000000000000000000000000",
282 => "000000000000000000000000",
283 => "000000000000000000000000",
284 => "000000000000000000000000",
285 => "000000000000000000000000",
286 => "000000000000000000000000",
287 => "000000000000000000000000",
288 => "000000000000000000000000",
289 => "000000000000000000000000",
290 => "000000000000000000000000",
291 => "000000000000000000000000",
292 => "000000000000000000000000",
293 => "000000000000000000000000",
294 => "000000000000000000000000",
295 => "000000000000000000000000",
296 => "000000000000000000000000",
297 => "000000000000000000000000",
298 => "000000000000000000000000",
299 => "000000000000000000000000",
300 => "000001110000011100000111",
301 => "111111111111111111111111",
302 => "111010011110100111101001",
303 => "101001001010010010100100",
304 => "010110010101100101011001",
305 => "001101100011011000110110",
306 => "111101001111010011110100",
307 => "100110101001101010011010",
308 => "111010101110101011101010",
309 => "100101101001011010010110",
310 => "001111100011111000111110",
311 => "111101111111011111110111",
312 => "111101001111010011110100",
313 => "001100110011001100110011",
314 => "111111001111110011111100",
315 => "110011001100110011001100",
316 => "010000010100000101000001",
317 => "111000111110001111100011",
318 => "100011101000111010001110",
319 => "111101011111010111110101",
320 => "111010111110101111101011",
321 => "001001010010010100100101",
322 => "100011011000110110001101",
323 => "110011111100111111001111",
324 => "100101011001010110010101",
325 => "111111101111111011111110",
326 => "011010100110101001101010",
327 => "000000000000000000000000",
328 => "000000000000000000000000",
329 => "000000000000000000000000",
330 => "100001111000011110000111",
331 => "111111111111111111111111",
332 => "001110110011101100111011",
333 => "000000000000000000000000",
334 => "001100110011001100110011",
335 => "010101100101011001010110",
336 => "001111110011111100111111",
337 => "111110101111101011111010",
338 => "111010001110100011101000",
339 => "001010000010100000101000",
340 => "110011001100110011001100",
341 => "111111111111111111111111",
342 => "011100000111000001110000",
343 => "101110001011100010111000",
344 => "111101001111010011110100",
345 => "011101000111010001110100",
346 => "111110011111100111111001",
347 => "111101111111011111110111",
348 => "111011101110111011101110",
349 => "101111001011110010111100",
350 => "111100111111001111110011",
351 => "111110111111101111111011",
352 => "010001010100010101000101",
353 => "000000000000000000000000",
354 => "000000000000000000000000",
355 => "000000000000000000000000",
356 => "000000000000000000000000",
357 => "000000000000000000000000",
358 => "000000000000000000000000",
359 => "000000000000000000000000",
360 => "000000000000000000000000",
361 => "000000000000000000000000",
362 => "000000000000000000000000",
363 => "000000000000000000000000",
364 => "000000000000000000000000",
365 => "000000000000000000000000",
366 => "000000000000000000000000",
367 => "000000000000000000000000",
368 => "000000000000000000000000",
369 => "000000000000000000000000",
370 => "000000000000000000000000",
371 => "000000000000000000000000",
372 => "000000000000000000000000",
373 => "000000000000000000000000",
374 => "000000000000000000000000",
375 => "000000000000000000000000",
376 => "000000000000000000000000",
377 => "000000000000000000000000",
378 => "000000000000000000000000",
379 => "000000000000000000000000",
380 => "000000000000000000000000",
381 => "000000000000000000000000",
382 => "000000000000000000000000",
383 => "000000000000000000000000",
384 => "000000000000000000000000",
385 => "000000000000000000000000",
386 => "000000000000000000000000",
387 => "000000000000000000000000",
388 => "000000000000000000000000",
389 => "000000000000000000000000",
390 => "000000000000000000000000",
391 => "000000000000000000000000",
392 => "000000000000000000000000",
393 => "000000000000000000000000",
394 => "000000000000000000000000",
395 => "000000000000000000000000",
396 => "000000000000000000000000",
397 => "000000000000000000000000",
398 => "000000000000000000000000",
399 => "000000000000000000000000",
400 => "000001110000011100000111",
401 => "111111111111111111111111",
402 => "111011111110111111101111",
403 => "101110011011100110111001",
404 => "011001100110011001100110",
405 => "100011111000111110001111",
406 => "111110111111101111111011",
407 => "101100011011000110110001",
408 => "110111101101111011011110",
409 => "110010111100101111001011",
410 => "000001110000011100000111",
411 => "101000011010000110100001",
412 => "111111111111111111111111",
413 => "100001111000011110000111",
414 => "111111011111110111111101",
415 => "010011100100111001001110",
416 => "000000000000000000000000",
417 => "000011010000110100001101",
418 => "101101001011010010110100",
419 => "111100001111000011110000",
420 => "010011110100111101001111",
421 => "000000000000000000000000",
422 => "000100010001000100010001",
423 => "010011110100111101001111",
424 => "100110101001101010011010",
425 => "111111001111110011111100",
426 => "100001111000011110000111",
427 => "000000000000000000000000",
428 => "000000000000000000000000",
429 => "000000000000000000000000",
430 => "100010111000101110001011",
431 => "111111111111111111111111",
432 => "010000010100000101000001",
433 => "000000000000000000000000",
434 => "000000000000000000000000",
435 => "000000000000000000000000",
436 => "000001100000011000000110",
437 => "110001011100010111000101",
438 => "111010001110100011101000",
439 => "000110010001100100011001",
440 => "010011100100111001001110",
441 => "111110111111101111111011",
442 => "101011001010110010101100",
443 => "111000001110000011100000",
444 => "101010101010101010101010",
445 => "000000100000001000000010",
446 => "110011111100111111001111",
447 => "111100111111001111110011",
448 => "001001010010010100100101",
449 => "001111000011110000111100",
450 => "100000111000001110000011",
451 => "111110111111101111111011",
452 => "010001010100010101000101",
453 => "000000000000000000000000",
454 => "000000000000000000000000",
455 => "000000000000000000000000",
456 => "000000000000000000000000",
457 => "000000000000000000000000",
458 => "000000000000000000000000",
459 => "000000000000000000000000",
460 => "000000000000000000000000",
461 => "000000000000000000000000",
462 => "000000000000000000000000",
463 => "000000000000000000000000",
464 => "000000000000000000000000",
465 => "000000000000000000000000",
466 => "000000000000000000000000",
467 => "000000000000000000000000",
468 => "000000000000000000000000",
469 => "000000000000000000000000",
470 => "000000000000000000000000",
471 => "000000000000000000000000",
472 => "000000000000000000000000",
473 => "000000000000000000000000",
474 => "000000000000000000000000",
475 => "000000000000000000000000",
476 => "000000000000000000000000",
477 => "000000000000000000000000",
478 => "000000000000000000000000",
479 => "000000000000000000000000",
480 => "000000000000000000000000",
481 => "000000000000000000000000",
482 => "000000000000000000000000",
483 => "000000000000000000000000",
484 => "000000000000000000000000",
485 => "000000000000000000000000",
486 => "000000000000000000000000",
487 => "000000000000000000000000",
488 => "000000000000000000000000",
489 => "000000000000000000000000",
490 => "000000000000000000000000",
491 => "000000000000000000000000",
492 => "000000000000000000000000",
493 => "000000000000000000000000",
494 => "000000000000000000000000",
495 => "000000000000000000000000",
496 => "000000000000000000000000",
497 => "000000000000000000000000",
498 => "000000000000000000000000",
499 => "000000000000000000000000",
500 => "000011010000110100001101",
501 => "111111111111111111111111",
502 => "110001011100010111000101",
503 => "000001000000010000000100",
504 => "000000000000000000000000",
505 => "100000111000001110000011",
506 => "111111101111111011111110",
507 => "100000001000000010000000",
508 => "010100110101001101010011",
509 => "100000011000000110000001",
510 => "000001010000010100000101",
511 => "001101000011010000110100",
512 => "111110011111100111111001",
513 => "111111001111110011111100",
514 => "110011001100110011001100",
515 => "000001000000010000000100",
516 => "000010100000101000001010",
517 => "101100101011001010110010",
518 => "111101011111010111110101",
519 => "011001100110011001100110",
520 => "101010001010100010101000",
521 => "001110110011101100111011",
522 => "110000001100000011000000",
523 => "110111101101111011011110",
524 => "011000100110001001100010",
525 => "111110011111100111111001",
526 => "100100111001001110010011",
527 => "000000100000001000000010",
528 => "000000000000000000000000",
529 => "000000000000000000000000",
530 => "010110000101100001011000",
531 => "111111101111111011111110",
532 => "110011001100110011001100",
533 => "001101010011010100110101",
534 => "001100000011000000110000",
535 => "011100000111000001110000",
536 => "000101010001010100010101",
537 => "110001011100010111000101",
538 => "111010001110100011101000",
539 => "000110010001100100011001",
540 => "000011000000110000001100",
541 => "110110101101101011011010",
542 => "111111101111111011111110",
543 => "111110101111101011111010",
544 => "001011110010111100101111",
545 => "000000000000000000000000",
546 => "110011111100111111001111",
547 => "111000101110001011100010",
548 => "000000010000000100000001",
549 => "000000000000000000000000",
550 => "100000111000001110000011",
551 => "111110111111101111111011",
552 => "010001010100010101000101",
553 => "000000000000000000000000",
554 => "000000000000000000000000",
555 => "000000000000000000000000",
556 => "000000000000000000000000",
557 => "000000000000000000000000",
558 => "000000000000000000000000",
559 => "000000000000000000000000",
560 => "000000000000000000000000",
561 => "000000000000000000000000",
562 => "000000000000000000000000",
563 => "000000000000000000000000",
564 => "000000000000000000000000",
565 => "000000000000000000000000",
566 => "000000000000000000000000",
567 => "000000000000000000000000",
568 => "000000000000000000000000",
569 => "000000000000000000000000",
570 => "000000000000000000000000",
571 => "000000000000000000000000",
572 => "000000000000000000000000",
573 => "000000000000000000000000",
574 => "000000000000000000000000",
575 => "000000000000000000000000",
576 => "000000000000000000000000",
577 => "000000000000000000000000",
578 => "000000000000000000000000",
579 => "000000000000000000000000",
580 => "000000000000000000000000",
581 => "000000000000000000000000",
582 => "000000000000000000000000",
583 => "000000000000000000000000",
584 => "000000000000000000000000",
585 => "000000000000000000000000",
586 => "000000000000000000000000",
587 => "000000000000000000000000",
588 => "000000000000000000000000",
589 => "000000000000000000000000",
590 => "000000000000000000000000",
591 => "000000000000000000000000",
592 => "000000000000000000000000",
593 => "000000000000000000000000",
594 => "000000000000000000000000",
595 => "000000000000000000000000",
596 => "000000000000000000000000",
597 => "000000000000000000000000",
598 => "000000000000000000000000",
599 => "000000000000000000000000",
600 => "100001001000010010000100",
601 => "111111111111111111111111",
602 => "111101001111010011110100",
603 => "010111110101111101011111",
604 => "000000000000000000000000",
605 => "001000110010001100100011",
606 => "110110111101101111011011",
607 => "111110011111100111111001",
608 => "111010001110100011101000",
609 => "101000011010000110100001",
610 => "000000110000001100000011",
611 => "000000100000001000000010",
612 => "101011101010111010101110",
613 => "111111111111111111111111",
614 => "010111000101110001011100",
615 => "000000000000000000000000",
616 => "010101100101011001010110",
617 => "111111111111111111111111",
618 => "111101011111010111110101",
619 => "110101001101010011010100",
620 => "111111001111110011111100",
621 => "010100000101000001010000",
622 => "110010101100101011001010",
623 => "111100011111000111110001",
624 => "110001011100010111000101",
625 => "111110101111101011111010",
626 => "111001001110010011100100",
627 => "000011100000111000001110",
628 => "000000000000000000000000",
629 => "000000000000000000000000",
630 => "000001100000011000000110",
631 => "101000011010000110100001",
632 => "111100111111001111110011",
633 => "111111111111111111111111",
634 => "111110101111101011111010",
635 => "110110001101100011011000",
636 => "010000000100000001000000",
637 => "111100011111000111110001",
638 => "111110011111100111111001",
639 => "011000110110001101100011",
640 => "000000000000000000000000",
641 => "011000000110000001100000",
642 => "111111101111111011111110",
643 => "101110011011100110111001",
644 => "000001000000010000000100",
645 => "001100110011001100110011",
646 => "111100101111001011110010",
647 => "111110011111100111111001",
648 => "011010000110100001101000",
649 => "000000000000000000000000",
650 => "111000001110000011100000",
651 => "111111101111111011111110",
652 => "101000111010001110100011",
653 => "000000000000000000000000",
654 => "000000000000000000000000",
655 => "000000000000000000000000",
656 => "000000000000000000000000",
657 => "000000000000000000000000",
658 => "000000000000000000000000",
659 => "000000000000000000000000",
660 => "000000000000000000000000",
661 => "000000000000000000000000",
662 => "000000000000000000000000",
663 => "000000000000000000000000",
664 => "000000000000000000000000",
665 => "000000000000000000000000",
666 => "000000000000000000000000",
667 => "000000000000000000000000",
668 => "000000000000000000000000",
669 => "000000000000000000000000",
670 => "000000000000000000000000",
671 => "000000000000000000000000",
672 => "000000000000000000000000",
673 => "000000000000000000000000",
674 => "000000000000000000000000",
675 => "000000000000000000000000",
676 => "000000000000000000000000",
677 => "000000000000000000000000",
678 => "000000000000000000000000",
679 => "000000000000000000000000",
680 => "000000000000000000000000",
681 => "000000000000000000000000",
682 => "000000000000000000000000",
683 => "000000000000000000000000",
684 => "000000000000000000000000",
685 => "000000000000000000000000",
686 => "000000000000000000000000",
687 => "000000000000000000000000",
688 => "000000000000000000000000",
689 => "000000000000000000000000",
690 => "000000000000000000000000",
691 => "000000000000000000000000",
692 => "000000000000000000000000",
693 => "000000000000000000000000",
694 => "000000000000000000000000",
695 => "000000000000000000000000",
696 => "000000000000000000000000",
697 => "000000000000000000000000",
698 => "000000000000000000000000",
699 => "000000000000000000000000",
700 => "001000110010001100100011",
701 => "001101110011011100110111",
702 => "001101110011011100110111",
703 => "000110010001100100011001",
704 => "000000000000000000000000",
705 => "000000000000000000000000",
706 => "000110000001100000011000",
707 => "001101100011011000110110",
708 => "001010110010101100101011",
709 => "000001010000010100000101",
710 => "000010110000101100001011",
711 => "001001110010011100100111",
712 => "100111001001110010011100",
713 => "110101011101010111010101",
714 => "000001100000011000000110",
715 => "000000000000000000000000",
716 => "000101000001010000010100",
717 => "001101110011011100110111",
718 => "001101110011011100110111",
719 => "001101110011011100110111",
720 => "001101110011011100110111",
721 => "000011110000111100001111",
722 => "000110010001100100011001",
723 => "001101100011011000110110",
724 => "001000000010000000100000",
725 => "001100010011000100110001",
726 => "001000000010000000100000",
727 => "000000010000000100000001",
728 => "000000000000000000000000",
729 => "000000000000000000000000",
730 => "000000000000000000000000",
731 => "000000110000001100000011",
732 => "001010000010100000101000",
733 => "001101110011011100110111",
734 => "001100010011000100110001",
735 => "000101000001010000010100",
736 => "000011010000110100001101",
737 => "001101110011011100110111",
738 => "001101110011011100110111",
739 => "000110110001101100011011",
740 => "000000000000000000000000",
741 => "000010100000101000001010",
742 => "001101100011011000110110",
743 => "000110110001101100011011",
744 => "000000000000000000000000",
745 => "000011110000111100001111",
746 => "001101110011011100110111",
747 => "001101110011011100110111",
748 => "000111100001111000011110",
749 => "000000000000000000000000",
750 => "001101110011011100110111",
751 => "001101110011011100110111",
752 => "001010100010101000101010",
753 => "000000000000000000000000",
754 => "000000000000000000000000",
755 => "000000000000000000000000",
756 => "000000000000000000000000",
757 => "000000000000000000000000",
758 => "000000000000000000000000",
759 => "000000000000000000000000",
760 => "000000000000000000000000",
761 => "000000000000000000000000",
762 => "000000000000000000000000",
763 => "000000000000000000000000",
764 => "000000000000000000000000",
765 => "000000000000000000000000",
766 => "000000000000000000000000",
767 => "000000000000000000000000",
768 => "000000000000000000000000",
769 => "000000000000000000000000",
770 => "000000000000000000000000",
771 => "000000000000000000000000",
772 => "000000000000000000000000",
773 => "000000000000000000000000",
774 => "000000000000000000000000",
775 => "000000000000000000000000",
776 => "000000000000000000000000",
777 => "000000000000000000000000",
778 => "000000000000000000000000",
779 => "000000000000000000000000",
780 => "000000000000000000000000",
781 => "000000000000000000000000",
782 => "000000000000000000000000",
783 => "000000000000000000000000",
784 => "000000000000000000000000",
785 => "000000000000000000000000",
786 => "000000000000000000000000",
787 => "000000000000000000000000",
788 => "000000000000000000000000",
789 => "000000000000000000000000",
790 => "000000000000000000000000",
791 => "000000000000000000000000",
792 => "000000000000000000000000",
793 => "000000000000000000000000",
794 => "000000000000000000000000",
795 => "000000000000000000000000",
796 => "000000000000000000000000",
797 => "000000000000000000000000",
798 => "000000000000000000000000",
799 => "000000000000000000000000",
800 => "000000000000000000000000",
801 => "000000000000000000000000",
802 => "000000000000000000000000",
803 => "000000000000000000000000",
804 => "000000000000000000000000",
805 => "000000000000000000000000",
806 => "000000000000000000000000",
807 => "000000000000000000000000",
808 => "000000000000000000000000",
809 => "000000000000000000000000",
810 => "001110110011101100111011",
811 => "111100111111001111110011",
812 => "111100011111000111110001",
813 => "010100010101000101010001",
814 => "000000000000000000000000",
815 => "000000000000000000000000",
816 => "000000000000000000000000",
817 => "000000000000000000000000",
818 => "000000000000000000000000",
819 => "000000000000000000000000",
820 => "000000000000000000000000",
821 => "000000000000000000000000",
822 => "000000000000000000000000",
823 => "000000000000000000000000",
824 => "000000000000000000000000",
825 => "000000000000000000000000",
826 => "000000000000000000000000",
827 => "000000000000000000000000",
828 => "000000000000000000000000",
829 => "000000000000000000000000",
830 => "000000000000000000000000",
831 => "000000000000000000000000",
832 => "000000000000000000000000",
833 => "000000000000000000000000",
834 => "000000000000000000000000",
835 => "000000000000000000000000",
836 => "000000000000000000000000",
837 => "000000000000000000000000",
838 => "000000000000000000000000",
839 => "000000000000000000000000",
840 => "000000000000000000000000",
841 => "000000000000000000000000",
842 => "000000000000000000000000",
843 => "000000000000000000000000",
844 => "000000000000000000000000",
845 => "000000000000000000000000",
846 => "000000000000000000000000",
847 => "000000000000000000000000",
848 => "000000000000000000000000",
849 => "000000000000000000000000",
850 => "000000000000000000000000",
851 => "000000000000000000000000",
852 => "000000000000000000000000",
853 => "000000000000000000000000",
854 => "000000000000000000000000",
855 => "000000000000000000000000",
856 => "000000000000000000000000",
857 => "000000000000000000000000",
858 => "000000000000000000000000",
859 => "000000000000000000000000",
860 => "000000000000000000000000",
861 => "000000000000000000000000",
862 => "000000000000000000000000",
863 => "000000000000000000000000",
864 => "000000000000000000000000",
865 => "000000000000000000000000",
866 => "000000000000000000000000",
867 => "000000000000000000000000",
868 => "000000000000000000000000",
869 => "000000000000000000000000",
870 => "000000000000000000000000",
871 => "000000000000000000000000",
872 => "000000000000000000000000",
873 => "000000000000000000000000",
874 => "000000000000000000000000",
875 => "000000000000000000000000",
876 => "000000000000000000000000",
877 => "000000000000000000000000",
878 => "000000000000000000000000",
879 => "000000000000000000000000",
880 => "000000000000000000000000",
881 => "000000000000000000000000",
882 => "000000000000000000000000",
883 => "000000000000000000000000",
884 => "000000000000000000000000",
885 => "000000000000000000000000",
886 => "000000000000000000000000",
887 => "000000000000000000000000",
888 => "000000000000000000000000",
889 => "000000000000000000000000",
890 => "000000000000000000000000",
891 => "000000000000000000000000",
892 => "000000000000000000000000",
893 => "000000000000000000000000",
894 => "000000000000000000000000",
895 => "000000000000000000000000",
896 => "000000000000000000000000",
897 => "000000000000000000000000",
898 => "000000000000000000000000",
899 => "000000000000000000000000",
900 => "000000000000000000000000",
901 => "000000000000000000000000",
902 => "000000000000000000000000",
903 => "000000000000000000000000",
904 => "000000000000000000000000",
905 => "000000000000000000000000",
906 => "000000000000000000000000",
907 => "000000000000000000000000",
908 => "000000000000000000000000",
909 => "000000000000000000000000",
910 => "000010010000100100001001",
911 => "001010000010100000101000",
912 => "001000000010000000100000",
913 => "000000000000000000000000",
914 => "000000000000000000000000",
915 => "000000000000000000000000",
916 => "000000000000000000000000",
917 => "000000000000000000000000",
918 => "000000000000000000000000",
919 => "000000000000000000000000",
920 => "000000000000000000000000",
921 => "000000000000000000000000",
922 => "000000000000000000000000",
923 => "000000000000000000000000",
924 => "000000000000000000000000",
925 => "000000000000000000000000",
926 => "000000000000000000000000",
927 => "000000000000000000000000",
928 => "000000000000000000000000",
929 => "000000000000000000000000",
930 => "000000000000000000000000",
931 => "000000000000000000000000",
932 => "000000000000000000000000",
933 => "000000000000000000000000",
934 => "000000000000000000000000",
935 => "000000000000000000000000",
936 => "000000000000000000000000",
937 => "000000000000000000000000",
938 => "000000000000000000000000",
939 => "000000000000000000000000",
940 => "000000000000000000000000",
941 => "000000000000000000000000",
942 => "000000000000000000000000",
943 => "000000000000000000000000",
944 => "000000000000000000000000",
945 => "000000000000000000000000",
946 => "000000000000000000000000",
947 => "000000000000000000000000",
948 => "000000000000000000000000",
949 => "000000000000000000000000",
950 => "000000000000000000000000",
951 => "000000000000000000000000",
952 => "000000000000000000000000",
953 => "000000000000000000000000",
954 => "000000000000000000000000",
955 => "000000000000000000000000",
956 => "000000000000000000000000",
957 => "000000000000000000000000",
958 => "000000000000000000000000",
959 => "000000000000000000000000",
960 => "000000000000000000000000",
961 => "000000000000000000000000",
962 => "000000000000000000000000",
963 => "000000000000000000000000",
964 => "000000000000000000000000",
965 => "000000000000000000000000",
966 => "000000000000000000000000",
967 => "000000000000000000000000",
968 => "000000000000000000000000",
969 => "000000000000000000000000",
970 => "000000000000000000000000",
971 => "000000000000000000000000",
972 => "000000000000000000000000",
973 => "000000000000000000000000",
974 => "000000000000000000000000",
975 => "000000000000000000000000",
976 => "000000000000000000000000",
977 => "000000000000000000000000",
978 => "000000000000000000000000",
979 => "000000000000000000000000",
980 => "000000000000000000000000",
981 => "000000000000000000000000",
982 => "000000000000000000000000",
983 => "000000000000000000000000",
984 => "000000000000000000000000",
985 => "000000000000000000000000",
986 => "000000000000000000000000",
987 => "000000000000000000000000",
988 => "000000000000000000000000",
989 => "000000000000000000000000",
990 => "000000000000000000000000",
991 => "000000000000000000000000",
992 => "000000000000000000000000",
993 => "000000000000000000000000",
994 => "000000000000000000000000",
995 => "000000000000000000000000",
996 => "000000000000000000000000",
997 => "000000000000000000000000",
998 => "000000000000000000000000",
999 => "000000000000000000000000",
1000 => "000000000000000000000000",
1001 => "000000000000000000000000",
1002 => "000000000000000000000000",
1003 => "000000000000000000000000",
1004 => "000000000000000000000000",
1005 => "000000000000000000000000",
1006 => "000000000000000000000000",
1007 => "000000000000000000000000",
1008 => "000000000000000000000000",
1009 => "000000000000000000000000",
1010 => "000000000000000000000000",
1011 => "000000000000000000000000",
1012 => "000000000000000000000000",
1013 => "000000000000000000000000",
1014 => "000000000000000000000000",
1015 => "000000000000000000000000",
1016 => "000000000000000000000000",
1017 => "000000000000000000000000",
1018 => "000000000000000000000000",
1019 => "000000000000000000000000",
1020 => "000000000000000000000000",
1021 => "000000000000000000000000",
1022 => "000000000000000000000000",
1023 => "000000000000000000000000",
1024 => "000000000000000000000000",
1025 => "000000000000000000000000",
1026 => "000000000000000000000000",
1027 => "000000000000000000000000",
1028 => "000000000000000000000000",
1029 => "000000000000000000000000",
1030 => "000000000000000000000000",
1031 => "000000000000000000000000",
1032 => "000000000000000000000000",
1033 => "000000000000000000000000",
1034 => "000000000000000000000000",
1035 => "000000000000000000000000",
1036 => "000000000000000000000000",
1037 => "000000000000000000000000",
1038 => "000000000000000000000000",
1039 => "000000000000000000000000",
1040 => "000000000000000000000000",
1041 => "000000000000000000000000",
1042 => "000000000000000000000000",
1043 => "000000000000000000000000",
1044 => "000000000000000000000000",
1045 => "000000000000000000000000",
1046 => "000000000000000000000000",
1047 => "000000000000000000000000",
1048 => "000000000000000000000000",
1049 => "000000000000000000000000",
1050 => "000000000000000000000000",
1051 => "000000000000000000000000",
1052 => "000000000000000000000000",
1053 => "000000000000000000000000",
1054 => "000000000000000000000000",
1055 => "000000000000000000000000",
1056 => "000000000000000000000000",
1057 => "000000000000000000000000",
1058 => "000000000000000000000000",
1059 => "000000000000000000000000",
1060 => "000000000000000000000000",
1061 => "000000000000000000000000",
1062 => "000000000000000000000000",
1063 => "000000000000000000000000",
1064 => "000000000000000000000000",
1065 => "000000000000000000000000",
1066 => "000000000000000000000000",
1067 => "000000000000000000000000",
1068 => "000000000000000000000000",
1069 => "000000000000000000000000",
1070 => "000000000000000000000000",
1071 => "000000000000000000000000",
1072 => "000000000000000000000000",
1073 => "000000000000000000000000",
1074 => "000000000000000000000000",
1075 => "000000000000000000000000",
1076 => "000000000000000000000000",
1077 => "000000000000000000000000",
1078 => "000000000000000000000000",
1079 => "000000000000000000000000",
1080 => "000000000000000000000000",
1081 => "000000000000000000000000",
1082 => "000000000000000000000000",
1083 => "000000000000000000000000",
1084 => "000000000000000000000000",
1085 => "000000000000000000000000",
1086 => "000000000000000000000000",
1087 => "000000000000000000000000",
1088 => "000000000000000000000000",
1089 => "000000000000000000000000",
1090 => "000000000000000000000000",
1091 => "000000000000000000000000",
1092 => "000000000000000000000000",
1093 => "000000000000000000000000",
1094 => "000000000000000000000000",
1095 => "000000000000000000000000",
1096 => "000000000000000000000000",
1097 => "000000000000000000000000",
1098 => "000000000000000000000000",
1099 => "000000000000000000000000",
1100 => "000000000000000000000000",
1101 => "000000000000000000000000",
1102 => "000000000000000000000000",
1103 => "000000000000000000000000",
1104 => "000000000000000000000000",
1105 => "000000000000000000000000",
1106 => "000000000000000000000000",
1107 => "000000000000000000000000",
1108 => "000000000000000000000000",
1109 => "000000000000000000000000",
1110 => "000000000000000000000000",
1111 => "000000000000000000000000",
1112 => "000000000000000000000000",
1113 => "000000000000000000000000",
1114 => "000000000000000000000000",
1115 => "000000000000000000000000",
1116 => "000000000000000000000000",
1117 => "000000000000000000000000",
1118 => "000000000000000000000000",
1119 => "000000000000000000000000",
1120 => "000000000000000000000000",
1121 => "000000000000000000000000",
1122 => "000000000000000000000000",
1123 => "000000000000000000000000",
1124 => "000000000000000000000000",
1125 => "000000000000000000000000",
1126 => "000000000000000000000000",
1127 => "000000000000000000000000",
1128 => "000000000000000000000000",
1129 => "000000000000000000000000",
1130 => "000000000000000000000000",
1131 => "000000000000000000000000",
1132 => "000000000000000000000000",
1133 => "000000000000000000000000",
1134 => "000000000000000000000000",
1135 => "000000000000000000000000",
1136 => "000000000000000000000000",
1137 => "000000000000000000000000",
1138 => "000000000000000000000000",
1139 => "000000010000000100000001",
1140 => "000011110000111100001111",
1141 => "000010100000101000001010",
1142 => "000000000000000000000000",
1143 => "000000000000000000000000",
1144 => "000000000000000000000000",
1145 => "000000000000000000000000",
1146 => "000000000000000000000000",
1147 => "000000000000000000000000",
1148 => "000000000000000000000000",
1149 => "000000000000000000000000",
1150 => "000000000000000000000000",
1151 => "000000000000000000000000",
1152 => "000000000000000000000000",
1153 => "000000000000000000000000",
1154 => "000000000000000000000000",
1155 => "000000000000000000000000",
1156 => "000000000000000000000000",
1157 => "000000000000000000000000",
1158 => "000000000000000000000000",
1159 => "000000000000000000000000",
1160 => "000000000000000000000000",
1161 => "000000000000000000000000",
1162 => "000000000000000000000000",
1163 => "000000000000000000000000",
1164 => "000000000000000000000000",
1165 => "000000000000000000000000",
1166 => "000000000000000000000000",
1167 => "000000000000000000000000",
1168 => "000000000000000000000000",
1169 => "000000000000000000000000",
1170 => "000000000000000000000000",
1171 => "000000000000000000000000",
1172 => "000000000000000000000000",
1173 => "000000000000000000000000",
1174 => "000000000000000000000000",
1175 => "000000000000000000000000",
1176 => "000000000000000000000000",
1177 => "000000000000000000000000",
1178 => "000000000000000000000000",
1179 => "000000000000000000000000",
1180 => "000000000000000000000000",
1181 => "000000000000000000000000",
1182 => "000000000000000000000000",
1183 => "000000000000000000000000",
1184 => "000000000000000000000000",
1185 => "000000010000000100000001",
1186 => "000100000001000000010000",
1187 => "000010100000101000001010",
1188 => "000000000000000000000000",
1189 => "000000000000000000000000",
1190 => "000000000000000000000000",
1191 => "000000000000000000000000",
1192 => "000000000000000000000000",
1193 => "000000000000000000000000",
1194 => "000000000000000000000000",
1195 => "000000000000000000000000",
1196 => "000000000000000000000000",
1197 => "000000000000000000000000",
1198 => "000000000000000000000000",
1199 => "000000000000000000000000",
1200 => "100100101001001010010010",
1201 => "111010001110100011101000",
1202 => "111010001110100011101000",
1203 => "111010001110100011101000",
1204 => "111010001110100011101000",
1205 => "010101110101011101010111",
1206 => "000000000000000000000000",
1207 => "000000000000000000000000",
1208 => "000000000000000000000000",
1209 => "000000000000000000000000",
1210 => "000000000000000000000000",
1211 => "000000000000000000000000",
1212 => "000000000000000000000000",
1213 => "000000000000000000000000",
1214 => "000000000000000000000000",
1215 => "000000000000000000000000",
1216 => "000000000000000000000000",
1217 => "000000000000000000000000",
1218 => "000000000000000000000000",
1219 => "000000000000000000000000",
1220 => "000000000000000000000000",
1221 => "000000000000000000000000",
1222 => "000000000000000000000000",
1223 => "000000000000000000000000",
1224 => "000000000000000000000000",
1225 => "000000000000000000000000",
1226 => "000000000000000000000000",
1227 => "011011010110110101101101",
1228 => "111010001110100011101000",
1229 => "111010001110100011101000",
1230 => "111010001110100011101000",
1231 => "111010001110100011101000",
1232 => "111010001110100011101000",
1233 => "101001111010011110100111",
1234 => "000000000000000000000000",
1235 => "000000000000000000000000",
1236 => "000000000000000000000000",
1237 => "000000000000000000000000",
1238 => "000000000000000000000000",
1239 => "101101111011011110110111",
1240 => "111011011110110111101101",
1241 => "100010101000101010001010",
1242 => "000000000000000000000000",
1243 => "000000000000000000000000",
1244 => "000000000000000000000000",
1245 => "000000000000000000000000",
1246 => "000000000000000000000000",
1247 => "000000000000000000000000",
1248 => "000000000000000000000000",
1249 => "000000000000000000000000",
1250 => "000000000000000000000000",
1251 => "000000000000000000000000",
1252 => "000000000000000000000000",
1253 => "000110110001101100011011",
1254 => "111010001110100011101000",
1255 => "111010001110100011101000",
1256 => "101110011011100110111001",
1257 => "110000101100001011000010",
1258 => "111010001110100011101000",
1259 => "110101011101010111010101",
1260 => "000011010000110100001101",
1261 => "000000000000000000000000",
1262 => "000000000000000000000000",
1263 => "000000000000000000000000",
1264 => "000000000000000000000000",
1265 => "000000000000000000000000",
1266 => "000000000000000000000000",
1267 => "000000000000000000000000",
1268 => "000000000000000000000000",
1269 => "000000000000000000000000",
1270 => "000000000000000000000000",
1271 => "000000000000000000000000",
1272 => "000000000000000000000000",
1273 => "000000000000000000000000",
1274 => "000000000000000000000000",
1275 => "000000000000000000000000",
1276 => "000000000000000000000000",
1277 => "000000000000000000000000",
1278 => "000000000000000000000000",
1279 => "000000000000000000000000",
1280 => "000000000000000000000000",
1281 => "000000000000000000000000",
1282 => "000000000000000000000000",
1283 => "000000000000000000000000",
1284 => "000001010000010100000101",
1285 => "101101111011011110110111",
1286 => "111011011110110111101101",
1287 => "100001011000010110000101",
1288 => "000000000000000000000000",
1289 => "000000000000000000000000",
1290 => "000000000000000000000000",
1291 => "000000000000000000000000",
1292 => "000000000000000000000000",
1293 => "000000000000000000000000",
1294 => "000000000000000000000000",
1295 => "000000000000000000000000",
1296 => "000000000000000000000000",
1297 => "000000000000000000000000",
1298 => "000000000000000000000000",
1299 => "000000000000000000000000",
1300 => "001010010010100100101001",
1301 => "111111111111111111111111",
1302 => "110110011101100111011001",
1303 => "011001000110010001100100",
1304 => "111010101110101011101010",
1305 => "011000000110000001100000",
1306 => "000000010000000100000001",
1307 => "000100010001000100010001",
1308 => "000100110001001100010011",
1309 => "010010000100100001001000",
1310 => "001100110011001100110011",
1311 => "000101000001010000010100",
1312 => "010011100100111001001110",
1313 => "001010100010101000101010",
1314 => "000000000000000000000000",
1315 => "010001100100011001000110",
1316 => "010100110101001101010011",
1317 => "001100000011000000110000",
1318 => "010010110100101101001011",
1319 => "000011100000111000001110",
1320 => "000100000001000000010000",
1321 => "010010110100101101001011",
1322 => "010001000100010001000100",
1323 => "000010110000101100001011",
1324 => "000000000000000000000000",
1325 => "000000000000000000000000",
1326 => "000000000000000000000000",
1327 => "011110000111100001111000",
1328 => "111001001110010011100100",
1329 => "100010111000101110001011",
1330 => "111111101111111011111110",
1331 => "101101011011010110110101",
1332 => "110000101100001011000010",
1333 => "101110001011100010111000",
1334 => "000111000001110000011100",
1335 => "010001110100011101000111",
1336 => "010100100101001001010010",
1337 => "001100100011001000110010",
1338 => "000000100000001000000010",
1339 => "001011110010111100101111",
1340 => "111100111111001111110011",
1341 => "100110101001101010011010",
1342 => "010001100100011001000110",
1343 => "001110110011101100111011",
1344 => "000000100000001000000010",
1345 => "000001100000011000000110",
1346 => "001101000011010000110100",
1347 => "010100110101001101010011",
1348 => "010010110100101101001011",
1349 => "000101000001010000010100",
1350 => "000000000000000000000000",
1351 => "000000000000000000000000",
1352 => "000000000000000000000000",
1353 => "000001100000011000000110",
1354 => "101001111010011110100111",
1355 => "111111111111111111111111",
1356 => "010101100101011001010110",
1357 => "101101011011010110110101",
1358 => "111101101111011011110110",
1359 => "011001010110010101100101",
1360 => "000000110000001100000011",
1361 => "000110100001101000011010",
1362 => "010001000100010001000100",
1363 => "010100110101001101010011",
1364 => "001101100011011000110110",
1365 => "000000000000000000000000",
1366 => "000111100001111000011110",
1367 => "010100110101001101010011",
1368 => "010011010100110101001101",
1369 => "001101010011010100110101",
1370 => "001100010011000100110001",
1371 => "001010100010101000101010",
1372 => "010011100100111001001110",
1373 => "010011110100111101001111",
1374 => "001000010010000100100001",
1375 => "000000000000000000000000",
1376 => "010010110100101101001011",
1377 => "010100110101001101010011",
1378 => "010010110100101101001011",
1379 => "001011100010111000101110",
1380 => "010100110101001101010011",
1381 => "001111110011111100111111",
1382 => "000000110000001100000011",
1383 => "000101000001010000010100",
1384 => "000010010000100100001001",
1385 => "001111100011111000111110",
1386 => "111111111111111111111111",
1387 => "100011101000111010001110",
1388 => "000001000000010000000100",
1389 => "001100100011001000110010",
1390 => "010100000101000001010000",
1391 => "010011010100110101001101",
1392 => "000101010001010100010101",
1393 => "000000000000000000000000",
1394 => "000001000000010000000100",
1395 => "000100110001001100010011",
1396 => "000101010001010100010101",
1397 => "010011110100111101001111",
1398 => "001010000010100000101000",
1399 => "000000000000000000000000",
1400 => "000001110000011100000111",
1401 => "111111111111111111111111",
1402 => "110110001101100011011000",
1403 => "010110100101101001011010",
1404 => "010010100100101001001010",
1405 => "000011110000111100001111",
1406 => "110011011100110111001101",
1407 => "111101001111010011110100",
1408 => "111010001110100011101000",
1409 => "111101111111011111110111",
1410 => "111101101111011011110110",
1411 => "110011001100110011001100",
1412 => "111111011111110111111101",
1413 => "111100001111000011110000",
1414 => "000011000000110000001100",
1415 => "110110001101100011011000",
1416 => "111111111111111111111111",
1417 => "111001001110010011100100",
1418 => "111101011111010111110101",
1419 => "001101010011010100110101",
1420 => "110011001100110011001100",
1421 => "110111011101110111011101",
1422 => "111001001110010011100100",
1423 => "101010111010101110101011",
1424 => "000000110000001100000011",
1425 => "000000000000000000000000",
1426 => "000000000000000000000000",
1427 => "000001110000011100000111",
1428 => "000010110000101100001011",
1429 => "010010000100100001001000",
1430 => "111111101111111011111110",
1431 => "100011011000110110001101",
1432 => "000010000000100000001000",
1433 => "000010110000101100001011",
1434 => "101000111010001110100011",
1435 => "111001101110011011100110",
1436 => "110100001101000011010000",
1437 => "111101011111010111110101",
1438 => "001111110011111100111111",
1439 => "001001000010010000100100",
1440 => "111100111111001111110011",
1441 => "111010101110101011101010",
1442 => "111101001111010011110100",
1443 => "111110111111101111111011",
1444 => "010000010100000101000001",
1445 => "001010100010101000101010",
1446 => "111101101111011011110110",
1447 => "101111101011111010111110",
1448 => "111101111111011111110111",
1449 => "110011101100111011001110",
1450 => "000000000000000000000000",
1451 => "000000000000000000000000",
1452 => "000000000000000000000000",
1453 => "000000000000000000000000",
1454 => "100011111000111110001111",
1455 => "111111111111111111111111",
1456 => "100100111001001110010011",
1457 => "111110101111101011111010",
1458 => "011111000111110001111100",
1459 => "000000100000001000000010",
1460 => "000000000000000000000000",
1461 => "100110111001101110011011",
1462 => "111010001110100011101000",
1463 => "110010101100101011001010",
1464 => "111110101111101011111010",
1465 => "010101110101011101010111",
1466 => "010111000101110001011100",
1467 => "111111111111111111111111",
1468 => "111010111110101111101011",
1469 => "111101101111011011110110",
1470 => "101000001010000010100000",
1471 => "110101101101011011010110",
1472 => "110100001101000011010000",
1473 => "111010001110100011101000",
1474 => "111001001110010011100100",
1475 => "000101000001010000010100",
1476 => "101110111011101110111011",
1477 => "111111111111111111111111",
1478 => "110100011101000111010001",
1479 => "011101000111010001110100",
1480 => "111111111111111111111111",
1481 => "100111111001111110011111",
1482 => "110011101100111011001110",
1483 => "111101001111010011110100",
1484 => "011011010110110101101101",
1485 => "001101000011010000110100",
1486 => "111111111111111111111111",
1487 => "100011101000111010001110",
1488 => "000111010001110100011101",
1489 => "111010111110101111101011",
1490 => "110000111100001111000011",
1491 => "111101001111010011110100",
1492 => "110011101100111011001110",
1493 => "000110100001101000011010",
1494 => "111001101110011011100110",
1495 => "111101001111010011110100",
1496 => "111001011110010111100101",
1497 => "111110111111101111111011",
1498 => "111011101110111011101110",
1499 => "000010110000101100001011",
1500 => "000001110000011100000111",
1501 => "111111111111111111111111",
1502 => "111110011111100111111001",
1503 => "111001011110010111100101",
1504 => "100111111001111110011111",
1505 => "000000000000000000000000",
1506 => "010001100100011001000110",
1507 => "111111111111111111111111",
1508 => "011110100111101001111010",
1509 => "100101011001010110010101",
1510 => "111111111111111111111111",
1511 => "010110010101100101011001",
1512 => "101101001011010010110100",
1513 => "111111111111111111111111",
1514 => "001001000010010000100100",
1515 => "010110110101101101011011",
1516 => "111111111111111111111111",
1517 => "100010001000100010001000",
1518 => "100010011000100110001001",
1519 => "011000110110001101100011",
1520 => "111111111111111111111111",
1521 => "100101001001010010010100",
1522 => "101010111010101110101011",
1523 => "111001101110011011100110",
1524 => "000101010001010100010101",
1525 => "000000000000000000000000",
1526 => "000000000000000000000000",
1527 => "000000000000000000000000",
1528 => "000000000000000000000000",
1529 => "010001110100011101000111",
1530 => "111111101111111011111110",
1531 => "100011011000110110001101",
1532 => "000000000000000000000000",
1533 => "000000000000000000000000",
1534 => "000010000000100000001000",
1535 => "001010110010101100101011",
1536 => "011110110111101101111011",
1537 => "111111111111111111111111",
1538 => "011000110110001101100011",
1539 => "001001000010010000100100",
1540 => "111100111111001111110011",
1541 => "101011101010111010101110",
1542 => "011000000110000001100000",
1543 => "111111111111111111111111",
1544 => "011111010111110101111101",
1545 => "000000100000001000000010",
1546 => "000101010001010100010101",
1547 => "001111000011110000111100",
1548 => "110100101101001011010010",
1549 => "111111111111111111111111",
1550 => "000000000000000000000000",
1551 => "000000000000000000000000",
1552 => "000000000000000000000000",
1553 => "000000000000000000000000",
1554 => "100011111000111110001111",
1555 => "111111111111111111111111",
1556 => "111101101111011011110110",
1557 => "111100111111001111110011",
1558 => "001100100011001000110010",
1559 => "000000000000000000000000",
1560 => "000000000000000000000000",
1561 => "000001100000011000000110",
1562 => "001010110010101100101011",
1563 => "011011110110111101101111",
1564 => "111111101111111011111110",
1565 => "100010001000100010001000",
1566 => "000001010000010100000101",
1567 => "110111111101111111011111",
1568 => "111010011110100111101001",
1569 => "010111010101110101011101",
1570 => "010111000101110001011100",
1571 => "000011010000110100001101",
1572 => "001101010011010100110101",
1573 => "101010111010101110101011",
1574 => "111111111111111111111111",
1575 => "000111110001111100011111",
1576 => "001000110010001100100011",
1577 => "111101011111010111110101",
1578 => "110101001101010011010100",
1579 => "011111110111111101111111",
1580 => "111101001111010011110100",
1581 => "000101010001010100010101",
1582 => "010111010101110101011101",
1583 => "111111111111111111111111",
1584 => "011100100111001001110010",
1585 => "001101000011010000110100",
1586 => "111111111111111111111111",
1587 => "100011101000111010001110",
1588 => "000000010000000100000001",
1589 => "000101000001010000010100",
1590 => "001111000011110000111100",
1591 => "110011011100110111001101",
1592 => "111010111110101111101011",
1593 => "000100000001000000010000",
1594 => "011111110111111101111111",
1595 => "111111111111111111111111",
1596 => "010111000101110001011100",
1597 => "101100011011000110110001",
1598 => "111111111111111111111111",
1599 => "000111110001111100011111",
1600 => "000001110000011100000111",
1601 => "111111111111111111111111",
1602 => "110001001100010011000100",
1603 => "000010000000100000001000",
1604 => "010100110101001101010011",
1605 => "001100110011001100110011",
1606 => "001101000011010000110100",
1607 => "111111111111111111111111",
1608 => "011010010110100101101001",
1609 => "100100101001001010010010",
1610 => "111111111111111111111111",
1611 => "001100100011001000110010",
1612 => "101001011010010110100101",
1613 => "111111111111111111111111",
1614 => "001001000010010000100100",
1615 => "010101100101011001010110",
1616 => "111111101111111011111110",
1617 => "010101100101011001010110",
1618 => "000000000000000000000000",
1619 => "010100100101001001010010",
1620 => "111111111111111111111111",
1621 => "101011101010111010101110",
1622 => "011100010111000101110001",
1623 => "100011001000110010001100",
1624 => "000100110001001100010011",
1625 => "000000000000000000000000",
1626 => "000000000000000000000000",
1627 => "000000000000000000000000",
1628 => "000000000000000000000000",
1629 => "010001110100011101000111",
1630 => "111111101111111011111110",
1631 => "100011011000110110001101",
1632 => "000000000000000000000000",
1633 => "000000100000001000000010",
1634 => "101100101011001010110010",
1635 => "110111111101111111011111",
1636 => "100011111000111110001111",
1637 => "111111111111111111111111",
1638 => "011000110110001101100011",
1639 => "001001000010010000100100",
1640 => "111100111111001111110011",
1641 => "100101001001010010010100",
1642 => "010010000100100001001000",
1643 => "111111111111111111111111",
1644 => "011111100111111001111110",
1645 => "010000000100000001000000",
1646 => "111100001111000011110000",
1647 => "101000111010001110100011",
1648 => "110010111100101111001011",
1649 => "111111111111111111111111",
1650 => "000000000000000000000000",
1651 => "000000000000000000000000",
1652 => "000000000000000000000000",
1653 => "000000000000000000000000",
1654 => "100011111000111110001111",
1655 => "111111111111111111111111",
1656 => "011011010110110101101101",
1657 => "111101001111010011110100",
1658 => "111000011110000111100001",
1659 => "000110110001101100011011",
1660 => "000001000000010000000100",
1661 => "101011101010111010101110",
1662 => "111000111110001111100011",
1663 => "100010111000101110001011",
1664 => "111111101111111011111110",
1665 => "100010001000100010001000",
1666 => "000000100000001000000010",
1667 => "110111101101111011011110",
1668 => "110010011100100111001001",
1669 => "000000000000000000000000",
1670 => "000110110001101100011011",
1671 => "110110011101100111011001",
1672 => "110000001100000011000000",
1673 => "101011011010110110101101",
1674 => "111111111111111111111111",
1675 => "000111110001111100011111",
1676 => "000000000000000000000000",
1677 => "101001101010011010100110",
1678 => "111111111111111111111111",
1679 => "111101111111011111110111",
1680 => "100101011001010110010101",
1681 => "000000000000000000000000",
1682 => "010110000101100001011000",
1683 => "111111111111111111111111",
1684 => "011100100111001001110010",
1685 => "001101000011010000110100",
1686 => "111111111111111111111111",
1687 => "100011101000111010001110",
1688 => "001100100011001000110010",
1689 => "111010101110101011101010",
1690 => "101010011010100110101001",
1691 => "110011001100110011001100",
1692 => "111010111110101111101011",
1693 => "000100000001000000010000",
1694 => "011110100111101001111010",
1695 => "111111111111111111111111",
1696 => "010010110100101101001011",
1697 => "101011111010111110101111",
1698 => "111111111111111111111111",
1699 => "000111110001111100011111",
1700 => "010111010101110101011101",
1701 => "111111111111111111111111",
1702 => "111011011110110111101101",
1703 => "101100101011001010110010",
1704 => "111100111111001111110011",
1705 => "100001101000011010000110",
1706 => "100001001000010010000100",
1707 => "111111111111111111111111",
1708 => "100111101001111010011110",
1709 => "100101111001011110010111",
1710 => "111111111111111111111111",
1711 => "011111010111110101111101",
1712 => "101001111010011110100111",
1713 => "111111111111111111111111",
1714 => "011000000110000001100000",
1715 => "100011001000110010001100",
1716 => "111111111111111111111111",
1717 => "100111011001110110011101",
1718 => "000000000000000000000000",
1719 => "000110000001100000011000",
1720 => "111001101110011011100110",
1721 => "111110001111100011111000",
1722 => "110110011101100111011001",
1723 => "110110011101100111011001",
1724 => "000100000001000000010000",
1725 => "000000000000000000000000",
1726 => "000000000000000000000000",
1727 => "000000000000000000000000",
1728 => "000011010000110100001101",
1729 => "101010101010101010101010",
1730 => "111111101111111011111110",
1731 => "110011001100110011001100",
1732 => "001001000010010000100100",
1733 => "000001010000010100000101",
1734 => "111110001111100011111000",
1735 => "110011101100111011001110",
1736 => "101011111010111110101111",
1737 => "111111111111111111111111",
1738 => "110010001100100011001000",
1739 => "100000101000001010000010",
1740 => "111110101111101011111010",
1741 => "110001111100011111000111",
1742 => "010101000101010001010100",
1743 => "111111111111111111111111",
1744 => "101010101010101010101010",
1745 => "011111100111111001111110",
1746 => "111111111111111111111111",
1747 => "100010101000101010001010",
1748 => "111100101111001011110010",
1749 => "111111111111111111111111",
1750 => "011110010111100101111001",
1751 => "000000000000000000000000",
1752 => "000000000000000000000000",
1753 => "000100000001000000010000",
1754 => "110011011100110111001101",
1755 => "111111111111111111111111",
1756 => "011000110110001101100011",
1757 => "110100001101000011010000",
1758 => "111111111111111111111111",
1759 => "110110101101101011011010",
1760 => "010001010100010101000101",
1761 => "111100111111001111110011",
1762 => "110101111101011111010111",
1763 => "101001011010010110100101",
1764 => "111111111111111111111111",
1765 => "111000011110000111100001",
1766 => "010001010100010101000101",
1767 => "111011001110110011101100",
1768 => "111001011110010111100101",
1769 => "001001100010011000100110",
1770 => "001111000011110000111100",
1771 => "111111111111111111111111",
1772 => "101010001010100010101000",
1773 => "110110001101100011011000",
1774 => "111111111111111111111111",
1775 => "101000111010001110100011",
1776 => "000001100000011000000110",
1777 => "001011010010110100101101",
1778 => "111110011111100111111001",
1779 => "111110011111100111111001",
1780 => "000111100001111000011110",
1781 => "000000000000000000000000",
1782 => "100011101000111010001110",
1783 => "111111111111111111111111",
1784 => "101010011010100110101001",
1785 => "011010010110100101101001",
1786 => "111111111111111111111111",
1787 => "101101101011011010110110",
1788 => "011101000111010001110100",
1789 => "111111111111111111111111",
1790 => "100100101001001010010010",
1791 => "111011011110110111101101",
1792 => "111111001111110011111100",
1793 => "100101101001011010010110",
1794 => "101011011010110110101101",
1795 => "111111111111111111111111",
1796 => "011111110111111101111111",
1797 => "101011111010111110101111",
1798 => "111111111111111111111111",
1799 => "011010010110100101101001",
1800 => "010110010101100101011001",
1801 => "100011101000111010001110",
1802 => "100011101000111010001110",
1803 => "100011101000111010001110",
1804 => "100011101000111010001110",
1805 => "010011100100111001001110",
1806 => "011110010111100101111001",
1807 => "100011101000111010001110",
1808 => "011110100111101001111010",
1809 => "010110000101100001011000",
1810 => "100011101000111010001110",
1811 => "011101000111010001110100",
1812 => "010111110101111101011111",
1813 => "100011101000111010001110",
1814 => "010111110101111101011111",
1815 => "011110010111100101111001",
1816 => "100011101000111010001110",
1817 => "100010011000100110001001",
1818 => "000000000000000000000000",
1819 => "000000000000000000000000",
1820 => "001001100010011000100110",
1821 => "100001001000010010000100",
1822 => "011111100111111001111110",
1823 => "000111010001110100011101",
1824 => "000000000000000000000000",
1825 => "000000000000000000000000",
1826 => "000000000000000000000000",
1827 => "000000000000000000000000",
1828 => "000011000000110000001100",
1829 => "100010111000101110001011",
1830 => "100011101000111010001110",
1831 => "100011101000111010001110",
1832 => "001000110010001100100011",
1833 => "000000010000000100000001",
1834 => "010010000100100001001000",
1835 => "100011001000110010001100",
1836 => "010100010101000101010001",
1837 => "011110110111101101111011",
1838 => "010011010100110101001101",
1839 => "011100110111001101110011",
1840 => "100011101000111010001110",
1841 => "100011101000111010001110",
1842 => "001110000011100000111000",
1843 => "100011101000111010001110",
1844 => "100000011000000110000001",
1845 => "000101010001010100010101",
1846 => "100000011000000110000001",
1847 => "011110100111101001111010",
1848 => "010100000101000001010000",
1849 => "100000001000000010000000",
1850 => "000111010001110100011101",
1851 => "000000000000000000000000",
1852 => "000000000000000000000000",
1853 => "000100010001000100010001",
1854 => "100011101000111010001110",
1855 => "100011101000111010001110",
1856 => "010010100100101001001010",
1857 => "011111010111110101111101",
1858 => "100011101000111010001110",
1859 => "100011101000111010001110",
1860 => "001100110011001100110011",
1861 => "010001010100010101000101",
1862 => "100011101000111010001110",
1863 => "010011100100111001001110",
1864 => "011111010111110101111101",
1865 => "010110000101100001011000",
1866 => "001101000011010000110100",
1867 => "100011101000111010001110",
1868 => "100011101000111010001110",
1869 => "001100110011001100110011",
1870 => "000001100000011000000110",
1871 => "011010010110100101101001",
1872 => "100001101000011010000110",
1873 => "010010000100100001001000",
1874 => "100000111000001110000011",
1875 => "001100100011001000110010",
1876 => "000000000000000000000000",
1877 => "000001010000010100000101",
1878 => "111000101110001011100010",
1879 => "101001111010011110100111",
1880 => "000000010000000100000001",
1881 => "000000000000000000000000",
1882 => "011110010111100101111001",
1883 => "100011101000111010001110",
1884 => "100010011000100110001001",
1885 => "011001000110010001100100",
1886 => "100011101000111010001110",
1887 => "100001001000010010000100",
1888 => "000111000001110000011100",
1889 => "011110010111100101111001",
1890 => "011111000111110001111100",
1891 => "010011000100110001001100",
1892 => "100000001000000010000000",
1893 => "001011010010110100101101",
1894 => "100001111000011110000111",
1895 => "100011101000111010001110",
1896 => "011100000111000001110000",
1897 => "011000110110001101100011",
1898 => "100011101000111010001110",
1899 => "011010010110100101101001",
1900 => "000000000000000000000000",
1901 => "000000000000000000000000",
1902 => "000000000000000000000000",
1903 => "000000000000000000000000",
1904 => "000000000000000000000000",
1905 => "000000000000000000000000",
1906 => "000000000000000000000000",
1907 => "000000000000000000000000",
1908 => "000000000000000000000000",
1909 => "000000000000000000000000",
1910 => "000000000000000000000000",
1911 => "000000000000000000000000",
1912 => "000000000000000000000000",
1913 => "000000000000000000000000",
1914 => "000000000000000000000000",
1915 => "000000000000000000000000",
1916 => "000000000000000000000000",
1917 => "000000000000000000000000",
1918 => "000000000000000000000000",
1919 => "000000000000000000000000",
1920 => "000000000000000000000000",
1921 => "000000000000000000000000",
1922 => "000000000000000000000000",
1923 => "000000000000000000000000",
1924 => "000000000000000000000000",
1925 => "000000000000000000000000",
1926 => "000000000000000000000000",
1927 => "000000000000000000000000",
1928 => "000000000000000000000000",
1929 => "000000000000000000000000",
1930 => "000000000000000000000000",
1931 => "000000000000000000000000",
1932 => "000000000000000000000000",
1933 => "000000000000000000000000",
1934 => "000000000000000000000000",
1935 => "000000000000000000000000",
1936 => "000000000000000000000000",
1937 => "000000000000000000000000",
1938 => "000000000000000000000000",
1939 => "000000000000000000000000",
1940 => "000000000000000000000000",
1941 => "000000000000000000000000",
1942 => "000000000000000000000000",
1943 => "000000000000000000000000",
1944 => "000000000000000000000000",
1945 => "000000000000000000000000",
1946 => "000000000000000000000000",
1947 => "000000000000000000000000",
1948 => "000000000000000000000000",
1949 => "000000000000000000000000",
1950 => "000000000000000000000000",
1951 => "000000000000000000000000",
1952 => "000000000000000000000000",
1953 => "000000000000000000000000",
1954 => "000000000000000000000000",
1955 => "000000000000000000000000",
1956 => "000000000000000000000000",
1957 => "000000000000000000000000",
1958 => "000000000000000000000000",
1959 => "000000000000000000000000",
1960 => "000000000000000000000000",
1961 => "000000000000000000000000",
1962 => "000000000000000000000000",
1963 => "000000000000000000000000",
1964 => "000000000000000000000000",
1965 => "000000000000000000000000",
1966 => "000000000000000000000000",
1967 => "000000000000000000000000",
1968 => "000000000000000000000000",
1969 => "000000000000000000000000",
1970 => "000000000000000000000000",
1971 => "000000000000000000000000",
1972 => "000000000000000000000000",
1973 => "000000000000000000000000",
1974 => "000000000000000000000000",
1975 => "000000000000000000000000",
1976 => "100100111001001110010011",
1977 => "110110011101100111011001",
1978 => "111101011111010111110101",
1979 => "001000110010001100100011",
1980 => "000000000000000000000000",
1981 => "000000000000000000000000",
1982 => "000000000000000000000000",
1983 => "000000000000000000000000",
1984 => "000000000000000000000000",
1985 => "000000000000000000000000",
1986 => "000000000000000000000000",
1987 => "000000000000000000000000",
1988 => "000000000000000000000000",
1989 => "000000000000000000000000",
1990 => "000000000000000000000000",
1991 => "000000000000000000000000",
1992 => "000000000000000000000000",
1993 => "000000000000000000000000",
1994 => "000000000000000000000000",
1995 => "000000000000000000000000",
1996 => "000000000000000000000000",
1997 => "000000000000000000000000",
1998 => "000000000000000000000000",
1999 => "000000000000000000000000",
2000 => "000000000000000000000000",
2001 => "000000000000000000000000",
2002 => "000000000000000000000000",
2003 => "000000000000000000000000",
2004 => "000000000000000000000000",
2005 => "000000000000000000000000",
2006 => "000000000000000000000000",
2007 => "000000000000000000000000",
2008 => "000000000000000000000000",
2009 => "000000000000000000000000",
2010 => "000000000000000000000000",
2011 => "000000000000000000000000",
2012 => "000000000000000000000000",
2013 => "000000000000000000000000",
2014 => "000000000000000000000000",
2015 => "000000000000000000000000",
2016 => "000000000000000000000000",
2017 => "000000000000000000000000",
2018 => "000000000000000000000000",
2019 => "000000000000000000000000",
2020 => "000000000000000000000000",
2021 => "000000000000000000000000",
2022 => "000000000000000000000000",
2023 => "000000000000000000000000",
2024 => "000000000000000000000000",
2025 => "000000000000000000000000",
2026 => "000000000000000000000000",
2027 => "000000000000000000000000",
2028 => "000000000000000000000000",
2029 => "000000000000000000000000",
2030 => "000000000000000000000000",
2031 => "000000000000000000000000",
2032 => "000000000000000000000000",
2033 => "000000000000000000000000",
2034 => "000000000000000000000000",
2035 => "000000000000000000000000",
2036 => "000000000000000000000000",
2037 => "000000000000000000000000",
2038 => "000000000000000000000000",
2039 => "000000000000000000000000",
2040 => "000000000000000000000000",
2041 => "000000000000000000000000",
2042 => "000000000000000000000000",
2043 => "000000000000000000000000",
2044 => "000000000000000000000000",
2045 => "000000000000000000000000",
2046 => "000000000000000000000000",
2047 => "000000000000000000000000",
2048 => "000000000000000000000000",
2049 => "000000000000000000000000",
2050 => "000000000000000000000000",
2051 => "000000000000000000000000",
2052 => "000000000000000000000000",
2053 => "000000000000000000000000",
2054 => "000000000000000000000000",
2055 => "000000000000000000000000",
2056 => "000000000000000000000000",
2057 => "000000000000000000000000",
2058 => "000000000000000000000000",
2059 => "000000000000000000000000",
2060 => "000000000000000000000000",
2061 => "000000000000000000000000",
2062 => "000000000000000000000000",
2063 => "000000000000000000000000",
2064 => "000000000000000000000000",
2065 => "000000000000000000000000",
2066 => "000000000000000000000000",
2067 => "000000000000000000000000",
2068 => "000000000000000000000000",
2069 => "000000000000000000000000",
2070 => "000000000000000000000000",
2071 => "000000000000000000000000",
2072 => "000000000000000000000000",
2073 => "000000000000000000000000",
2074 => "000000000000000000000000",
2075 => "000000000000000000000000",
2076 => "010011000100110001001100",
2077 => "100000101000001010000010",
2078 => "001111010011110100111101",
2079 => "000000000000000000000000",
2080 => "000000000000000000000000",
2081 => "000000000000000000000000",
2082 => "000000000000000000000000",
2083 => "000000000000000000000000",
2084 => "000000000000000000000000",
2085 => "000000000000000000000000",
2086 => "000000000000000000000000",
2087 => "000000000000000000000000",
2088 => "000000000000000000000000",
2089 => "000000000000000000000000",
2090 => "000000000000000000000000",
2091 => "000000000000000000000000",
2092 => "000000000000000000000000",
2093 => "000000000000000000000000",
2094 => "000000000000000000000000",
2095 => "000000000000000000000000",
2096 => "000000000000000000000000",
2097 => "000000000000000000000000",
2098 => "000000000000000000000000",
2099 => "000000000000000000000000",
2100 => "000000000000000000000000",
2101 => "000000000000000000000000",
2102 => "000000000000000000000000",
2103 => "000000000000000000000000",
2104 => "000000000000000000000000",
2105 => "000000000000000000000000",
2106 => "000000000000000000000000",
2107 => "000000000000000000000000",
2108 => "000000000000000000000000",
2109 => "000000000000000000000000",
2110 => "000000000000000000000000",
2111 => "000000000000000000000000",
2112 => "000000000000000000000000",
2113 => "000000000000000000000000",
2114 => "000000000000000000000000",
2115 => "000000000000000000000000",
2116 => "000000000000000000000000",
2117 => "000000000000000000000000",
2118 => "000000000000000000000000",
2119 => "000000000000000000000000",
2120 => "000000000000000000000000",
2121 => "000000000000000000000000",
2122 => "000000000000000000000000",
2123 => "000000000000000000000000",
2124 => "000000000000000000000000",
2125 => "000000000000000000000000",
2126 => "000000000000000000000000",
2127 => "000000000000000000000000",
2128 => "000000000000000000000000",
2129 => "000000000000000000000000",
2130 => "000000000000000000000000",
2131 => "000000000000000000000000",
2132 => "000000000000000000000000",
2133 => "000000000000000000000000",
2134 => "000000000000000000000000",
2135 => "000000000000000000000000",
2136 => "000000000000000000000000",
2137 => "000000000000000000000000",
2138 => "000000000000000000000000",
2139 => "000000000000000000000000",
2140 => "000000000000000000000000",
2141 => "000000000000000000000000",
2142 => "000000000000000000000000",
2143 => "000000000000000000000000",
2144 => "000000000000000000000000",
2145 => "000000000000000000000000",
2146 => "000000000000000000000000",
2147 => "000000000000000000000000",
2148 => "000000000000000000000000",
2149 => "000000000000000000000000",
2150 => "000000000000000000000000",
2151 => "000000000000000000000000",
2152 => "000000000000000000000000",
2153 => "000000000000000000000000",
2154 => "000000000000000000000000",
2155 => "000000000000000000000000",
2156 => "000000000000000000000000",
2157 => "000000000000000000000000",
2158 => "000000000000000000000000",
2159 => "000000000000000000000000",
2160 => "000000000000000000000000",
2161 => "000000000000000000000000",
2162 => "000000000000000000000000",
2163 => "000000000000000000000000",
2164 => "000000000000000000000000",
2165 => "000000000000000000000000",
2166 => "000000000000000000000000",
2167 => "000000000000000000000000",
2168 => "000000000000000000000000",
2169 => "000000000000000000000000",
2170 => "000000000000000000000000",
2171 => "000000000000000000000000",
2172 => "000000000000000000000000",
2173 => "000000000000000000000000",
2174 => "000000000000000000000000",
2175 => "000000000000000000000000",
2176 => "000000000000000000000000",
2177 => "000000000000000000000000",
2178 => "000000000000000000000000",
2179 => "000000000000000000000000",
2180 => "000000000000000000000000",
2181 => "000000000000000000000000",
2182 => "000000000000000000000000",
2183 => "000000000000000000000000",
2184 => "000000000000000000000000",
2185 => "000000000000000000000000",
2186 => "000000000000000000000000",
2187 => "000000000000000000000000",
2188 => "000000000000000000000000",
2189 => "000000000000000000000000",
2190 => "000000000000000000000000",
2191 => "000000000000000000000000",
2192 => "000000000000000000000000",
2193 => "000000000000000000000000",
2194 => "000000000000000000000000",
2195 => "000000000000000000000000",
2196 => "000000000000000000000000",
2197 => "000000000000000000000000",
2198 => "000000000000000000000000",
2199 => "000000000000000000000000",
2200 => "000000000000000000000000",
2201 => "000000000000000000000000",
2202 => "000000000000000000000000",
2203 => "000000000000000000000000",
2204 => "000000000000000000000000",
2205 => "000000000000000000000000",
2206 => "000000000000000000000000",
2207 => "000000010000000100000001",
2208 => "000000110000001100000011",
2209 => "000000010000000100000001",
2210 => "000001010000010100000101",
2211 => "000010110000101100001011",
2212 => "000000110000001100000011",
2213 => "000011000000110000001100",
2214 => "000011000000110000001100",
2215 => "000001100000011000000110",
2216 => "000000000000000000000000",
2217 => "000000000000000000000000",
2218 => "000000000000000000000000",
2219 => "000000000000000000000000",
2220 => "000000000000000000000000",
2221 => "000000000000000000000000",
2222 => "000000000000000000000000",
2223 => "000000000000000000000000",
2224 => "000000000000000000000000",
2225 => "000000000000000000000000",
2226 => "000000000000000000000000",
2227 => "000000000000000000000000",
2228 => "000000000000000000000000",
2229 => "000000100000001000000010",
2230 => "000000110000001100000011",
2231 => "000000010000000100000001",
2232 => "000000000000000000000000",
2233 => "000000000000000000000000",
2234 => "000000000000000000000000",
2235 => "000000000000000000000000",
2236 => "000000000000000000000000",
2237 => "000000000000000000000000",
2238 => "000000000000000000000000",
2239 => "000000000000000000000000",
2240 => "000000000000000000000000",
2241 => "000000000000000000000000",
2242 => "000000000000000000000000",
2243 => "000000000000000000000000",
2244 => "000000000000000000000000",
2245 => "000000000000000000000000",
2246 => "000000000000000000000000",
2247 => "000000000000000000000000",
2248 => "000000000000000000000000",
2249 => "000000000000000000000000",
2250 => "000000000000000000000000",
2251 => "000000000000000000000000",
2252 => "000000010000000100000001",
2253 => "000010100000101000001010",
2254 => "000010000000100000001000",
2255 => "000000000000000000000000",
2256 => "000000000000000000000000",
2257 => "000000000000000000000000",
2258 => "000000000000000000000000",
2259 => "000000000000000000000000",
2260 => "000000000000000000000000",
2261 => "000000000000000000000000",
2262 => "000000000000000000000000",
2263 => "000000000000000000000000",
2264 => "000000000000000000000000",
2265 => "000000000000000000000000",
2266 => "000000000000000000000000",
2267 => "000000000000000000000000",
2268 => "000000000000000000000000",
2269 => "000000000000000000000000",
2270 => "000000000000000000000000",
2271 => "000000000000000000000000",
2272 => "000000000000000000000000",
2273 => "000000000000000000000000",
2274 => "000000000000000000000000",
2275 => "000000000000000000000000",
2276 => "000000000000000000000000",
2277 => "000000000000000000000000",
2278 => "000000000000000000000000",
2279 => "000000000000000000000000",
2280 => "000000000000000000000000",
2281 => "000000000000000000000000",
2282 => "000000000000000000000000",
2283 => "000000000000000000000000",
2284 => "000000000000000000000000",
2285 => "000000000000000000000000",
2286 => "000000000000000000000000",
2287 => "000000000000000000000000",
2288 => "000000000000000000000000",
2289 => "000000000000000000000000",
2290 => "000000000000000000000000",
2291 => "000000000000000000000000",
2292 => "000000000000000000000000",
2293 => "000000000000000000000000",
2294 => "000000000000000000000000",
2295 => "000000000000000000000000",
2296 => "000000000000000000000000",
2297 => "000000000000000000000000",
2298 => "000000000000000000000000",
2299 => "000000000000000000000000",
2300 => "000000000000000000000000",
2301 => "000000100000001000000010",
2302 => "011010010110100101101001",
2303 => "100110011001100110011001",
2304 => "001101000011010000110100",
2305 => "000000000000000000000000",
2306 => "000101110001011100010111",
2307 => "100110001001100010011000",
2308 => "101100011011000110110001",
2309 => "001011010010110100101101",
2310 => "100110011001100110011001",
2311 => "111110111111101111111011",
2312 => "010110100101101001011010",
2313 => "111011011110110111101101",
2314 => "111111111111111111111111",
2315 => "100010001000100010001000",
2316 => "000000000000000000000000",
2317 => "000000000000000000000000",
2318 => "000000000000000000000000",
2319 => "000000000000000000000000",
2320 => "000000000000000000000000",
2321 => "000000000000000000000000",
2322 => "000000000000000000000000",
2323 => "000000000000000000000000",
2324 => "000000000000000000000000",
2325 => "000000000000000000000000",
2326 => "000000000000000000000000",
2327 => "000000000000000000000000",
2328 => "001010000010100000101000",
2329 => "101001011010010110100101",
2330 => "101100111011001110110011",
2331 => "000111010001110100011101",
2332 => "000000000000000000000000",
2333 => "000000000000000000000000",
2334 => "000000000000000000000000",
2335 => "000000000000000000000000",
2336 => "000000000000000000000000",
2337 => "000000010000000100000001",
2338 => "001101100011011000110110",
2339 => "100100011001000110010001",
2340 => "100101011001010110010101",
2341 => "011001100110011001100110",
2342 => "000010000000100000001000",
2343 => "000000000000000000000000",
2344 => "000000000000000000000000",
2345 => "000000000000000000000000",
2346 => "000000000000000000000000",
2347 => "000000000000000000000000",
2348 => "000000000000000000000000",
2349 => "000000000000000000000000",
2350 => "000000000000000000000000",
2351 => "000000000000000000000000",
2352 => "001000110010001100100011",
2353 => "111100001111000011110000",
2354 => "110011011100110111001101",
2355 => "000010100000101000001010",
2356 => "000000000000000000000000",
2357 => "000000000000000000000000",
2358 => "000000000000000000000000",
2359 => "000000000000000000000000",
2360 => "000000000000000000000000",
2361 => "000000000000000000000000",
2362 => "000000000000000000000000",
2363 => "000000000000000000000000",
2364 => "000000000000000000000000",
2365 => "000000000000000000000000",
2366 => "000000000000000000000000",
2367 => "000000000000000000000000",
2368 => "000000000000000000000000",
2369 => "000000000000000000000000",
2370 => "000000000000000000000000",
2371 => "000000000000000000000000",
2372 => "000000000000000000000000",
2373 => "000000000000000000000000",
2374 => "000000000000000000000000",
2375 => "000000000000000000000000",
2376 => "000000000000000000000000",
2377 => "000000000000000000000000",
2378 => "000000000000000000000000",
2379 => "000000000000000000000000",
2380 => "000000000000000000000000",
2381 => "000000000000000000000000",
2382 => "000000000000000000000000",
2383 => "000000000000000000000000",
2384 => "000000000000000000000000",
2385 => "000000000000000000000000",
2386 => "000000000000000000000000",
2387 => "000000000000000000000000",
2388 => "000000000000000000000000",
2389 => "000000000000000000000000",
2390 => "000000000000000000000000",
2391 => "000000000000000000000000",
2392 => "000000000000000000000000",
2393 => "000000000000000000000000",
2394 => "000000000000000000000000",
2395 => "000000000000000000000000",
2396 => "000000000000000000000000",
2397 => "000000000000000000000000",
2398 => "000000000000000000000000",
2399 => "000000000000000000000000",
2400 => "000000000000000000000000",
2401 => "000011010000110100001101",
2402 => "111001011110010111100101",
2403 => "111111101111111011111110",
2404 => "101010001010100010101000",
2405 => "000000010000000100000001",
2406 => "000011010000110100001101",
2407 => "101010111010101110101011",
2408 => "111111111111111111111111",
2409 => "001111110011111100111111",
2410 => "001011000010110000101100",
2411 => "010111100101111001011110",
2412 => "000110000001100000011000",
2413 => "010010110100101101001011",
2414 => "111111101111111011111110",
2415 => "100010111000101110001011",
2416 => "000101010001010100010101",
2417 => "000100000001000000010000",
2418 => "000000000000000000000000",
2419 => "000000000000000000000000",
2420 => "000010010000100100001001",
2421 => "000101110001011100010111",
2422 => "000100000001000000010000",
2423 => "000000010000000100000001",
2424 => "000011000000110000001100",
2425 => "000110000001100000011000",
2426 => "000111000001110000011100",
2427 => "000100100001001000010010",
2428 => "001000110010001100100011",
2429 => "110001101100011011000110",
2430 => "111111111111111111111111",
2431 => "001010110010101100101011",
2432 => "000110000001100000011000",
2433 => "000110000001100000011000",
2434 => "000010000000100000001000",
2435 => "000000000000000000000000",
2436 => "000000000000000000000000",
2437 => "000111100001111000011110",
2438 => "111100001111000011110000",
2439 => "101111011011110110111101",
2440 => "100111001001110010011100",
2441 => "111111111111111111111111",
2442 => "000111010001110100011101",
2443 => "000000000000000000000000",
2444 => "000010110000101100001011",
2445 => "000110000001100000011000",
2446 => "000011110000111100001111",
2447 => "000000000000000000000000",
2448 => "000011100000111000001110",
2449 => "000110000001100000011000",
2450 => "000110000001100000011000",
2451 => "000100110001001100010011",
2452 => "000011110000111100001111",
2453 => "010101110101011101010111",
2454 => "010001100100011001000110",
2455 => "000000100000001000000010",
2456 => "000000100000001000000010",
2457 => "000001010000010100000101",
2458 => "000010110000101100001011",
2459 => "000101100001011000010110",
2460 => "000001100000011000000110",
2461 => "000000000000000000000000",
2462 => "000000000000000000000000",
2463 => "000000000000000000000000",
2464 => "000000000000000000000000",
2465 => "000000000000000000000000",
2466 => "000000000000000000000000",
2467 => "000000000000000000000000",
2468 => "000000000000000000000000",
2469 => "000000000000000000000000",
2470 => "000000000000000000000000",
2471 => "000000000000000000000000",
2472 => "000000000000000000000000",
2473 => "000000000000000000000000",
2474 => "000000000000000000000000",
2475 => "000000000000000000000000",
2476 => "000000000000000000000000",
2477 => "000000000000000000000000",
2478 => "000000000000000000000000",
2479 => "000000000000000000000000",
2480 => "000000000000000000000000",
2481 => "000000000000000000000000",
2482 => "000000000000000000000000",
2483 => "000000000000000000000000",
2484 => "000000000000000000000000",
2485 => "000000000000000000000000",
2486 => "000000000000000000000000",
2487 => "000000000000000000000000",
2488 => "000000000000000000000000",
2489 => "000000000000000000000000",
2490 => "000000000000000000000000",
2491 => "000000000000000000000000",
2492 => "000000000000000000000000",
2493 => "000000000000000000000000",
2494 => "000000000000000000000000",
2495 => "000000000000000000000000",
2496 => "000000000000000000000000",
2497 => "000000000000000000000000",
2498 => "000000000000000000000000",
2499 => "000000000000000000000000",
2500 => "000000000000000000000000",
2501 => "010010110100101101001011",
2502 => "111100011111000111110001",
2503 => "110001111100011111000111",
2504 => "111001111110011111100111",
2505 => "000101100001011000010110",
2506 => "000000000000000000000000",
2507 => "100000111000001110000011",
2508 => "111111111111111111111111",
2509 => "001111110011111100111111",
2510 => "101000111010001110100011",
2511 => "110000001100000011000000",
2512 => "010110010101100101011001",
2513 => "010010110100101101001011",
2514 => "111111101111111011111110",
2515 => "111000011110000111100001",
2516 => "111100111111001111110011",
2517 => "111000011110000111100001",
2518 => "001001110010011100100111",
2519 => "000100110001001100010011",
2520 => "101111111011111110111111",
2521 => "111010111110101111101011",
2522 => "110111111101111111011111",
2523 => "010001010100010101000101",
2524 => "100001011000010110000101",
2525 => "111111111111111111111111",
2526 => "110111001101110011011100",
2527 => "111010011110100111101001",
2528 => "011110010111100101111001",
2529 => "101001111010011110100111",
2530 => "111111111111111111111111",
2531 => "011100000111000001110000",
2532 => "111111111111111111111111",
2533 => "111101111111011111110111",
2534 => "010010010100100101001001",
2535 => "000000000000000000000000",
2536 => "000000000000000000000000",
2537 => "001010100010101000101010",
2538 => "111110001111100011111000",
2539 => "101110011011100110111001",
2540 => "001101000011010000110100",
2541 => "010101000101010001010100",
2542 => "000010010000100100001001",
2543 => "001000000010000000100000",
2544 => "110011011100110111001101",
2545 => "111010111110101111101011",
2546 => "111000001110000011100000",
2547 => "001110010011100100111001",
2548 => "100101011001010110010101",
2549 => "111111111111111111111111",
2550 => "110011001100110011001100",
2551 => "111011101110111011101110",
2552 => "100110101001101010011010",
2553 => "101110101011101010111010",
2554 => "101010111010101110101011",
2555 => "001010010010100100101001",
2556 => "101101011011010110110101",
2557 => "101111001011110010111100",
2558 => "110011001100110011001100",
2559 => "111110101111101011111010",
2560 => "100101001001010010010100",
2561 => "000000100000001000000010",
2562 => "000000000000000000000000",
2563 => "000000000000000000000000",
2564 => "000000000000000000000000",
2565 => "000000000000000000000000",
2566 => "000000000000000000000000",
2567 => "000000000000000000000000",
2568 => "000000000000000000000000",
2569 => "000000000000000000000000",
2570 => "000000000000000000000000",
2571 => "000000000000000000000000",
2572 => "000000000000000000000000",
2573 => "000000000000000000000000",
2574 => "000000000000000000000000",
2575 => "000000000000000000000000",
2576 => "000000000000000000000000",
2577 => "000000000000000000000000",
2578 => "000000000000000000000000",
2579 => "000000000000000000000000",
2580 => "000000000000000000000000",
2581 => "000000000000000000000000",
2582 => "000000000000000000000000",
2583 => "000000000000000000000000",
2584 => "000000000000000000000000",
2585 => "000000000000000000000000",
2586 => "000000000000000000000000",
2587 => "000000000000000000000000",
2588 => "000000000000000000000000",
2589 => "000000000000000000000000",
2590 => "000000000000000000000000",
2591 => "000000000000000000000000",
2592 => "000000000000000000000000",
2593 => "000000000000000000000000",
2594 => "000000000000000000000000",
2595 => "000000000000000000000000",
2596 => "000000000000000000000000",
2597 => "000000000000000000000000",
2598 => "000000000000000000000000",
2599 => "000000000000000000000000",
2600 => "000000100000001000000010",
2601 => "101010101010101010101010",
2602 => "110000011100000111000001",
2603 => "011010000110100001101000",
2604 => "111111011111110111111101",
2605 => "010011100100111001001110",
2606 => "000000000000000000000000",
2607 => "100000111000001110000011",
2608 => "111111111111111111111111",
2609 => "001111110011111100111111",
2610 => "011111010111110101111101",
2611 => "111111111111111111111111",
2612 => "011101010111010101110101",
2613 => "010010110100101101001011",
2614 => "111111101111111011111110",
2615 => "101011011010110110101101",
2616 => "100000111000001110000011",
2617 => "111111111111111111111111",
2618 => "011110010111100101111001",
2619 => "011110010111100101111001",
2620 => "111101101111011011110110",
2621 => "010101110101011101010111",
2622 => "110101011101010111010101",
2623 => "101111101011111010111110",
2624 => "001111000011110000111100",
2625 => "111100111111001111110011",
2626 => "110110111101101111011011",
2627 => "101001101010011010100110",
2628 => "011010000110100001101000",
2629 => "101001111010011110100111",
2630 => "111111111111111111111111",
2631 => "100011001000110010001100",
2632 => "111111101111111011111110",
2633 => "011010100110101001101010",
2634 => "000000000000000000000000",
2635 => "000000000000000000000000",
2636 => "000000000000000000000000",
2637 => "000000110000001100000011",
2638 => "011100010111000101110001",
2639 => "111011011110110111101101",
2640 => "111100001111000011110000",
2641 => "100100001001000010010000",
2642 => "000010100000101000001010",
2643 => "100100111001001110010011",
2644 => "111101011111010111110101",
2645 => "010000010100000101000001",
2646 => "111000101110001011100010",
2647 => "101010001010100010101000",
2648 => "001111100011111000111110",
2649 => "111111111111111111111111",
2650 => "110101111101011111010111",
2651 => "101010111010101110101011",
2652 => "011100100111001001110010",
2653 => "110111111101111111011111",
2654 => "111000111110001111100011",
2655 => "000110110001101100011011",
2656 => "110110111101101111011011",
2657 => "111110001111100011111000",
2658 => "010111000101110001011100",
2659 => "111100001111000011110000",
2660 => "110100111101001111010011",
2661 => "000001110000011100000111",
2662 => "000000000000000000000000",
2663 => "000000000000000000000000",
2664 => "000000000000000000000000",
2665 => "000000000000000000000000",
2666 => "000000000000000000000000",
2667 => "000000000000000000000000",
2668 => "000000000000000000000000",
2669 => "000000000000000000000000",
2670 => "000000000000000000000000",
2671 => "000000000000000000000000",
2672 => "000000000000000000000000",
2673 => "000000000000000000000000",
2674 => "000000000000000000000000",
2675 => "000000000000000000000000",
2676 => "000000000000000000000000",
2677 => "000000000000000000000000",
2678 => "000000000000000000000000",
2679 => "000000000000000000000000",
2680 => "000000000000000000000000",
2681 => "000000000000000000000000",
2682 => "000000000000000000000000",
2683 => "000000000000000000000000",
2684 => "000000000000000000000000",
2685 => "000000000000000000000000",
2686 => "000000000000000000000000",
2687 => "000000000000000000000000",
2688 => "000000000000000000000000",
2689 => "000000000000000000000000",
2690 => "000000000000000000000000",
2691 => "000000000000000000000000",
2692 => "000000000000000000000000",
2693 => "000000000000000000000000",
2694 => "000000000000000000000000",
2695 => "000000000000000000000000",
2696 => "000000000000000000000000",
2697 => "000000000000000000000000",
2698 => "000000000000000000000000",
2699 => "000000000000000000000000",
2700 => "000100110001001100010011",
2701 => "111011111110111111101111",
2702 => "111011111110111111101111",
2703 => "111010101110101011101010",
2704 => "111111001111110011111100",
2705 => "101101001011010010110100",
2706 => "000000100000001000000010",
2707 => "100000111000001110000011",
2708 => "111111111111111111111111",
2709 => "001111110011111100111111",
2710 => "010100100101001001010010",
2711 => "111111111111111111111111",
2712 => "011101010111010101110101",
2713 => "010010110100101101001011",
2714 => "111111101111111011111110",
2715 => "011010110110101101101011",
2716 => "010000010100000101000001",
2717 => "111111111111111111111111",
2718 => "100000111000001110000011",
2719 => "101000001010000010100000",
2720 => "111111001111110011111100",
2721 => "101111011011110110111101",
2722 => "101011011010110110101101",
2723 => "101000111010001110100011",
2724 => "001000110010001100100011",
2725 => "111011101110111011101110",
2726 => "101101011011010110110101",
2727 => "000000010000000100000001",
2728 => "000000000000000000000000",
2729 => "101001111010011110100111",
2730 => "111111111111111111111111",
2731 => "111100011111000111110001",
2732 => "111111011111110111111101",
2733 => "001101100011011000110110",
2734 => "000000000000000000000000",
2735 => "000000000000000000000000",
2736 => "000000000000000000000000",
2737 => "000010110000101100001011",
2738 => "001010000010100000101000",
2739 => "001011100010111000101110",
2740 => "101111001011110010111100",
2741 => "111111101111111011111110",
2742 => "010100100101001001010010",
2743 => "101110111011101110111011",
2744 => "111111001111110011111100",
2745 => "101100111011001110110011",
2746 => "101011011010110110101101",
2747 => "100101011001010110010101",
2748 => "000111000001110000011100",
2749 => "111111111111111111111111",
2750 => "100111001001110010011100",
2751 => "000000000000000000000000",
2752 => "000010100000101000001010",
2753 => "110100101101001011010010",
2754 => "111000111110001111100011",
2755 => "000011100000111000001110",
2756 => "110011001100110011001100",
2757 => "111011101110111011101110",
2758 => "001010000010100000101000",
2759 => "111010111110101111101011",
2760 => "110100111101001111010011",
2761 => "000001110000011100000111",
2762 => "000000000000000000000000",
2763 => "000000000000000000000000",
2764 => "000000000000000000000000",
2765 => "000000000000000000000000",
2766 => "000000000000000000000000",
2767 => "000000000000000000000000",
2768 => "000000000000000000000000",
2769 => "000000000000000000000000",
2770 => "000000000000000000000000",
2771 => "000000000000000000000000",
2772 => "000000000000000000000000",
2773 => "000000000000000000000000",
2774 => "000000000000000000000000",
2775 => "000000000000000000000000",
2776 => "000000000000000000000000",
2777 => "000000000000000000000000",
2778 => "000000000000000000000000",
2779 => "000000000000000000000000",
2780 => "000000000000000000000000",
2781 => "000000000000000000000000",
2782 => "000000000000000000000000",
2783 => "000000000000000000000000",
2784 => "000000000000000000000000",
2785 => "000000000000000000000000",
2786 => "000000000000000000000000",
2787 => "000000000000000000000000",
2788 => "000000000000000000000000",
2789 => "000000000000000000000000",
2790 => "000000000000000000000000",
2791 => "000000000000000000000000",
2792 => "000000000000000000000000",
2793 => "000000000000000000000000",
2794 => "000000000000000000000000",
2795 => "000000000000000000000000",
2796 => "000000000000000000000000",
2797 => "000000000000000000000000",
2798 => "000000000000000000000000",
2799 => "000000000000000000000000",
2800 => "011110110111101101111011",
2801 => "111110111111101111111011",
2802 => "011011000110110001101100",
2803 => "001101100011011000110110",
2804 => "111001001110010011100100",
2805 => "111011101110111011101110",
2806 => "010010010100100101001001",
2807 => "100101101001011010010110",
2808 => "111111111111111111111111",
2809 => "010110000101100001011000",
2810 => "011011110110111101101111",
2811 => "111111111111111111111111",
2812 => "100010101000101010001010",
2813 => "010011000100110001001100",
2814 => "111111101111111011111110",
2815 => "110011011100110111001101",
2816 => "101111001011110010111100",
2817 => "111110101111101011111010",
2818 => "010000110100001101000011",
2819 => "010110100101101001011010",
2820 => "111110111111101111111011",
2821 => "110010101100101011001010",
2822 => "101001101010011010100110",
2823 => "101100101011001010110010",
2824 => "001100000011000000110000",
2825 => "111100011111000111110001",
2826 => "110001001100010011000100",
2827 => "000010110000101100001011",
2828 => "000010000000100000001000",
2829 => "101111001011110010111100",
2830 => "111111111111111111111111",
2831 => "011100000111000001110000",
2832 => "111111111111111111111111",
2833 => "110100111101001111010011",
2834 => "000110100001101000011010",
2835 => "000000000000000000000000",
2836 => "000000000000000000000000",
2837 => "010001010100010101000101",
2838 => "111110111111101111111011",
2839 => "011001110110011101100111",
2840 => "100100001001000010010000",
2841 => "111110101111101011111010",
2842 => "010001010100010101000101",
2843 => "011100100111001001110010",
2844 => "111111101111111011111110",
2845 => "110000001100000011000000",
2846 => "101011001010110010101100",
2847 => "100110011001100110011001",
2848 => "001100100011001000110010",
2849 => "111111111111111111111111",
2850 => "101011111010111110101111",
2851 => "000010010000100100001001",
2852 => "000110000001100000011000",
2853 => "110110111101101111011011",
2854 => "111010001110100011101000",
2855 => "001001100010011000100110",
2856 => "110101101101011011010110",
2857 => "111100101111001011110010",
2858 => "001111100011111000111110",
2859 => "111010111110101111101011",
2860 => "111000011110000111100001",
2861 => "000111010001110100011101",
2862 => "000000000000000000000000",
2863 => "000000000000000000000000",
2864 => "000000000000000000000000",
2865 => "000000000000000000000000",
2866 => "000000000000000000000000",
2867 => "000000000000000000000000",
2868 => "000000000000000000000000",
2869 => "000000000000000000000000",
2870 => "000000000000000000000000",
2871 => "000000000000000000000000",
2872 => "000000000000000000000000",
2873 => "000000000000000000000000",
2874 => "000000000000000000000000",
2875 => "000000000000000000000000",
2876 => "000000000000000000000000",
2877 => "000000000000000000000000",
2878 => "000000000000000000000000",
2879 => "000000000000000000000000",
2880 => "000000000000000000000000",
2881 => "000000000000000000000000",
2882 => "000000000000000000000000",
2883 => "000000000000000000000000",
2884 => "000000000000000000000000",
2885 => "000000000000000000000000",
2886 => "000000000000000000000000",
2887 => "000000000000000000000000",
2888 => "000000000000000000000000",
2889 => "000000000000000000000000",
2890 => "000000000000000000000000",
2891 => "000000000000000000000000",
2892 => "000000000000000000000000",
2893 => "000000000000000000000000",
2894 => "000000000000000000000000",
2895 => "000000000000000000000000",
2896 => "000000000000000000000000",
2897 => "000000000000000000000000",
2898 => "000000000000000000000000",
2899 => "000000000000000000000000",
2900 => "101011101010111010101110",
2901 => "110010101100101011001010",
2902 => "011111100111111001111110",
2903 => "001100100011001000110010",
2904 => "110010101100101011001010",
2905 => "110010101100101011001010",
2906 => "100100101001001010010010",
2907 => "101110001011100010111000",
2908 => "110010101100101011001010",
2909 => "100111011001110110011101",
2910 => "101111101011111010111110",
2911 => "110010101100101011001010",
2912 => "101101001011010010110100",
2913 => "001111110011111100111111",
2914 => "110000001100000011000000",
2915 => "011101110111011101110111",
2916 => "110010011100100111001001",
2917 => "011010100110101001101010",
2918 => "000000110000001100000011",
2919 => "000001110000011100000111",
2920 => "011101000111010001110100",
2921 => "110001001100010011000100",
2922 => "101001001010010010100100",
2923 => "001011000010110000101100",
2924 => "011010010110100101101001",
2925 => "110010101100101011001010",
2926 => "110010101100101011001010",
2927 => "001010110010101100101011",
2928 => "001000100010001000100010",
2929 => "110001101100011011000110",
2930 => "110010101100101011001010",
2931 => "001100010011000100110001",
2932 => "110010011100100111001001",
2933 => "110010101100101011001010",
2934 => "010110100101101001011010",
2935 => "000000000000000000000000",
2936 => "000000000000000000000000",
2937 => "000111100001111000011110",
2938 => "100111001001110010011100",
2939 => "110001111100011111000111",
2940 => "110000001100000011000000",
2941 => "010110110101101101011011",
2942 => "000000110000001100000011",
2943 => "000010010000100100001001",
2944 => "100000111000001110000011",
2945 => "110010001100100011001000",
2946 => "100111011001110110011101",
2947 => "001001010010010100100101",
2948 => "011101100111011001110110",
2949 => "110010101100101011001010",
2950 => "110001101100011011000110",
2951 => "001010000010100000101000",
2952 => "010001000100010001000100",
2953 => "110010101100101011001010",
2954 => "110010101100101011001010",
2955 => "011011110110111101101111",
2956 => "110010101100101011001010",
2957 => "110010101100101011001010",
2958 => "011111110111111101111111",
2959 => "101110101011101010111010",
2960 => "110010101100101011001010",
2961 => "011000100110001001100010",
2962 => "000000000000000000000000",
2963 => "000000000000000000000000",
2964 => "000000000000000000000000",
2965 => "000000000000000000000000",
2966 => "000000000000000000000000",
2967 => "000000000000000000000000",
2968 => "000000000000000000000000",
2969 => "000000000000000000000000",
2970 => "000000000000000000000000",
2971 => "000000000000000000000000",
2972 => "000000000000000000000000",
2973 => "000000000000000000000000",
2974 => "000000000000000000000000",
2975 => "000000000000000000000000",
2976 => "000000000000000000000000",
2977 => "000000000000000000000000",
2978 => "000000000000000000000000",
2979 => "000000000000000000000000",
2980 => "000000000000000000000000",
2981 => "000000000000000000000000",
2982 => "000000000000000000000000",
2983 => "000000000000000000000000",
2984 => "000000000000000000000000",
2985 => "000000000000000000000000",
2986 => "000000000000000000000000",
2987 => "000000000000000000000000",
2988 => "000000000000000000000000",
2989 => "000000000000000000000000",
2990 => "000000000000000000000000",
2991 => "000000000000000000000000",
2992 => "000000000000000000000000",
2993 => "000000000000000000000000",
2994 => "000000000000000000000000",
2995 => "000000000000000000000000",
2996 => "000000000000000000000000",
2997 => "000000000000000000000000",
2998 => "000000000000000000000000",
2999 => "000000000000000000000000",
3000 => "000000000000000000000000",
3001 => "000000000000000000000000",
3002 => "000000000000000000000000",
3003 => "000000000000000000000000",
3004 => "000000000000000000000000",
3005 => "000000000000000000000000",
3006 => "000000000000000000000000",
3007 => "000000000000000000000000",
3008 => "000000000000000000000000",
3009 => "000000000000000000000000",
3010 => "000000000000000000000000",
3011 => "000000000000000000000000",
3012 => "000000000000000000000000",
3013 => "000000000000000000000000",
3014 => "000000000000000000000000",
3015 => "000000000000000000000000",
3016 => "000000000000000000000000",
3017 => "000000000000000000000000",
3018 => "000000000000000000000000",
3019 => "000000000000000000000000",
3020 => "000000000000000000000000",
3021 => "000000000000000000000000",
3022 => "000000000000000000000000",
3023 => "000000000000000000000000",
3024 => "000000000000000000000000",
3025 => "000000000000000000000000",
3026 => "000000000000000000000000",
3027 => "000000000000000000000000",
3028 => "000000000000000000000000",
3029 => "000000000000000000000000",
3030 => "000000000000000000000000",
3031 => "000000000000000000000000",
3032 => "000000000000000000000000",
3033 => "000000000000000000000000",
3034 => "000000000000000000000000",
3035 => "000000000000000000000000",
3036 => "000000000000000000000000",
3037 => "000000000000000000000000",
3038 => "000000000000000000000000",
3039 => "000000000000000000000000",
3040 => "000000000000000000000000",
3041 => "000000000000000000000000",
3042 => "000000000000000000000000",
3043 => "000000000000000000000000",
3044 => "000000000000000000000000",
3045 => "000000000000000000000000",
3046 => "000000000000000000000000",
3047 => "000000000000000000000000",
3048 => "000000000000000000000000",
3049 => "000000000000000000000000",
3050 => "000000000000000000000000",
3051 => "000000000000000000000000",
3052 => "000000000000000000000000",
3053 => "000000000000000000000000",
3054 => "000000000000000000000000",
3055 => "000000000000000000000000",
3056 => "000000000000000000000000",
3057 => "000000000000000000000000",
3058 => "000000000000000000000000",
3059 => "000000000000000000000000",
3060 => "000000000000000000000000",
3061 => "000000000000000000000000",
3062 => "000000000000000000000000",
3063 => "000000000000000000000000",
3064 => "000000000000000000000000",
3065 => "000000000000000000000000",
3066 => "000000000000000000000000",
3067 => "000000000000000000000000",
3068 => "000000000000000000000000",
3069 => "000000000000000000000000",
3070 => "000000000000000000000000",
3071 => "000000000000000000000000",
3072 => "000000000000000000000000",
3073 => "000000000000000000000000",
3074 => "000000000000000000000000",
3075 => "000000000000000000000000",
3076 => "000000000000000000000000",
3077 => "000000000000000000000000",
3078 => "000000000000000000000000",
3079 => "000000000000000000000000",
3080 => "000000000000000000000000",
3081 => "000000000000000000000000",
3082 => "000000000000000000000000",
3083 => "000000000000000000000000",
3084 => "000000000000000000000000",
3085 => "000000000000000000000000",
3086 => "000000000000000000000000",
3087 => "000000000000000000000000",
3088 => "000000000000000000000000",
3089 => "000000000000000000000000",
3090 => "000000000000000000000000",
3091 => "000000000000000000000000",
3092 => "000000000000000000000000",
3093 => "000000000000000000000000",
3094 => "000000000000000000000000",
3095 => "000000000000000000000000",
3096 => "000000000000000000000000",
3097 => "000000000000000000000000",
3098 => "000000000000000000000000",
3099 => "000000000000000000000000",
3100 => "000000000000000000000000",
3101 => "000000000000000000000000",
3102 => "000000000000000000000000",
3103 => "000000000000000000000000",
3104 => "000000000000000000000000",
3105 => "000000000000000000000000",
3106 => "000000000000000000000000",
3107 => "000000000000000000000000",
3108 => "000000000000000000000000",
3109 => "000000000000000000000000",
3110 => "000000000000000000000000",
3111 => "000000000000000000000000",
3112 => "000000000000000000000000",
3113 => "000000000000000000000000",
3114 => "000000000000000000000000",
3115 => "000000000000000000000000",
3116 => "000000000000000000000000",
3117 => "000000000000000000000000",
3118 => "000000000000000000000000",
3119 => "000000000000000000000000",
3120 => "000000000000000000000000",
3121 => "000000000000000000000000",
3122 => "000000000000000000000000",
3123 => "000000000000000000000000",
3124 => "000000000000000000000000",
3125 => "000000000000000000000000",
3126 => "000000000000000000000000",
3127 => "000000000000000000000000",
3128 => "000000000000000000000000",
3129 => "000000000000000000000000",
3130 => "000000000000000000000000",
3131 => "000000000000000000000000",
3132 => "000000000000000000000000",
3133 => "000000000000000000000000",
3134 => "000000000000000000000000",
3135 => "000000000000000000000000",
3136 => "000000000000000000000000",
3137 => "000000000000000000000000",
3138 => "000000000000000000000000",
3139 => "000000000000000000000000",
3140 => "000000000000000000000000",
3141 => "000000000000000000000000",
3142 => "000000000000000000000000",
3143 => "000000000000000000000000",
3144 => "000000000000000000000000",
3145 => "000000000000000000000000",
3146 => "000000000000000000000000",
3147 => "000000000000000000000000",
3148 => "000000000000000000000000",
3149 => "000000000000000000000000",
3150 => "000000000000000000000000",
3151 => "000000000000000000000000",
3152 => "000000000000000000000000",
3153 => "000000000000000000000000",
3154 => "000000000000000000000000",
3155 => "000000000000000000000000",
3156 => "000000000000000000000000",
3157 => "000000000000000000000000",
3158 => "000000000000000000000000",
3159 => "000000000000000000000000",
3160 => "000000000000000000000000",
3161 => "000000000000000000000000",
3162 => "000000000000000000000000",
3163 => "000000000000000000000000",
3164 => "000000000000000000000000",
3165 => "000000000000000000000000",
3166 => "000000000000000000000000",
3167 => "000000000000000000000000",
3168 => "000000000000000000000000",
3169 => "000000000000000000000000",
3170 => "000000000000000000000000",
3171 => "000000000000000000000000",
3172 => "000000000000000000000000",
3173 => "000000000000000000000000",
3174 => "000000000000000000000000",
3175 => "000000000000000000000000",
3176 => "000000000000000000000000",
3177 => "000000000000000000000000",
3178 => "000000000000000000000000",
3179 => "000000000000000000000000",
3180 => "000000000000000000000000",
3181 => "000000000000000000000000",
3182 => "000000000000000000000000",
3183 => "000000000000000000000000",
3184 => "000000000000000000000000",
3185 => "000000000000000000000000",
3186 => "000000000000000000000000",
3187 => "000000000000000000000000",
3188 => "000000000000000000000000",
3189 => "000000000000000000000000",
3190 => "000000000000000000000000",
3191 => "000000000000000000000000",
3192 => "000000000000000000000000",
3193 => "000000000000000000000000",
3194 => "000000000000000000000000",
3195 => "000000000000000000000000",
3196 => "000000000000000000000000",
3197 => "000000000000000000000000",
3198 => "000000000000000000000000",
3199 => "000000000000000000000000",
3200 => "000000000000000000000000",
3201 => "000000000000000000000000",
3202 => "000000000000000000000000",
3203 => "000000000000000000000000",
3204 => "000000000000000000000000",
3205 => "000000000000000000000000",
3206 => "000000000000000000000000",
3207 => "000000000000000000000000",
3208 => "000000000000000000000000",
3209 => "000000000000000000000000",
3210 => "000000000000000000000000",
3211 => "000000000000000000000000",
3212 => "000000000000000000000000",
3213 => "000000000000000000000000",
3214 => "000000000000000000000000",
3215 => "000000000000000000000000",
3216 => "000000000000000000000000",
3217 => "000000000000000000000000",
3218 => "000000000000000000000000",
3219 => "000000000000000000000000",
3220 => "000000000000000000000000",
3221 => "000000000000000000000000",
3222 => "000000000000000000000000",
3223 => "000000000000000000000000",
3224 => "000000000000000000000000",
3225 => "000000000000000000000000",
3226 => "000000000000000000000000",
3227 => "000000000000000000000000",
3228 => "000000000000000000000000",
3229 => "000000000000000000000000",
3230 => "000000000000000000000000",
3231 => "000000000000000000000000",
3232 => "000000000000000000000000",
3233 => "000000000000000000000000",
3234 => "000000000000000000000000",
3235 => "000000000000000000000000",
3236 => "000000000000000000000000",
3237 => "000000000000000000000000",
3238 => "000000000000000000000000",
3239 => "000000000000000000000000",
3240 => "000000000000000000000000",
3241 => "000000000000000000000000",
3242 => "000000000000000000000000",
3243 => "000000000000000000000000",
3244 => "000000000000000000000000",
3245 => "000000000000000000000000",
3246 => "000000000000000000000000",
3247 => "000000000000000000000000",
3248 => "000000000000000000000000",
3249 => "000000000000000000000000",
3250 => "000000000000000000000000",
3251 => "000000000000000000000000",
3252 => "000000000000000000000000",
3253 => "000000000000000000000000",
3254 => "000000000000000000000000",
3255 => "000000000000000000000000",
3256 => "000000000000000000000000",
3257 => "000000000000000000000000",
3258 => "000000000000000000000000",
3259 => "000000000000000000000000",
3260 => "000000000000000000000000",
3261 => "000000000000000000000000",
3262 => "000000000000000000000000",
3263 => "000000000000000000000000",
3264 => "000000000000000000000000",
3265 => "000000000000000000000000",
3266 => "000000000000000000000000",
3267 => "000000000000000000000000",
3268 => "000000000000000000000000",
3269 => "000000000000000000000000",
3270 => "000000000000000000000000",
3271 => "000000000000000000000000",
3272 => "000000000000000000000000",
3273 => "000000000000000000000000",
3274 => "000000000000000000000000",
3275 => "000000000000000000000000",
3276 => "000000000000000000000000",
3277 => "000000000000000000000000",
3278 => "000000000000000000000000",
3279 => "000000000000000000000000",
3280 => "000000000000000000000000",
3281 => "000000000000000000000000",
3282 => "000000000000000000000000",
3283 => "000000000000000000000000",
3284 => "000000000000000000000000",
3285 => "000000000000000000000000",
3286 => "000000000000000000000000",
3287 => "000000000000000000000000",
3288 => "000000000000000000000000",
3289 => "000000000000000000000000",
3290 => "000000000000000000000000",
3291 => "000000000000000000000000",
3292 => "000000000000000000000000",
3293 => "000000000000000000000000",
3294 => "000000000000000000000000",
3295 => "000000000000000000000000",
3296 => "000000000000000000000000",
3297 => "000000000000000000000000",
3298 => "000000000000000000000000",
3299 => "000000000000000000000000",
3300 => "000000000000000000000000",
3301 => "000000000000000000000000",
3302 => "000000000000000000000000",
3303 => "000000000000000000000000",
3304 => "000000000000000000000000",
3305 => "000000000000000000000000",
3306 => "000000000000000000000000",
3307 => "000000000000000000000000",
3308 => "000000000000000000000000",
3309 => "000000000000000000000000",
3310 => "000000000000000000000000",
3311 => "000000000000000000000000",
3312 => "000000000000000000000000",
3313 => "000000000000000000000000",
3314 => "000000000000000000000000",
3315 => "000000000000000000000000",
3316 => "000000000000000000000000",
3317 => "000000000000000000000000",
3318 => "000000000000000000000000",
3319 => "000000000000000000000000",
3320 => "000000000000000000000000",
3321 => "000000000000000000000000",
3322 => "000000000000000000000000",
3323 => "000000000000000000000000",
3324 => "000000000000000000000000",
3325 => "000000000000000000000000",
3326 => "000000000000000000000000",
3327 => "000000000000000000000000",
3328 => "000000000000000000000000",
3329 => "000000000000000000000000",
3330 => "000000000000000000000000",
3331 => "000000000000000000000000",
3332 => "000000000000000000000000",
3333 => "000000000000000000000000",
3334 => "000000000000000000000000",
3335 => "000000000000000000000000",
3336 => "000000000000000000000000",
3337 => "000000000000000000000000",
3338 => "000000000000000000000000",
3339 => "000000000000000000000000",
3340 => "000000000000000000000000",
3341 => "000000000000000000000000",
3342 => "000000000000000000000000",
3343 => "000000000000000000000000",
3344 => "000000000000000000000000",
3345 => "000000000000000000000000",
3346 => "000000000000000000000000",
3347 => "000000000000000000000000",
3348 => "000000000000000000000000",
3349 => "000000000000000000000000",
3350 => "000000000000000000000000",
3351 => "000000000000000000000000",
3352 => "000000000000000000000000",
3353 => "000000000000000000000000",
3354 => "000000000000000000000000",
3355 => "000000000000000000000000",
3356 => "000000000000000000000000",
3357 => "000000000000000000000000",
3358 => "000000000000000000000000",
3359 => "000000000000000000000000",
3360 => "000000000000000000000000",
3361 => "000000000000000000000000",
3362 => "000000000000000000000000",
3363 => "000000000000000000000000",
3364 => "000000000000000000000000",
3365 => "000000000000000000000000",
3366 => "000000000000000000000000",
3367 => "000000000000000000000000",
3368 => "000000000000000000000000",
3369 => "000000000000000000000000",
3370 => "000000000000000000000000",
3371 => "000000000000000000000000",
3372 => "000000000000000000000000",
3373 => "000000000000000000000000",
3374 => "000000000000000000000000",
3375 => "000000000000000000000000",
3376 => "000000000000000000000000",
3377 => "000000000000000000000000",
3378 => "000000000000000000000000",
3379 => "000000000000000000000000",
3380 => "000000000000000000000000",
3381 => "000000000000000000000000",
3382 => "000000000000000000000000",
3383 => "000000000000000000000000",
3384 => "000000000000000000000000",
3385 => "000000000000000000000000",
3386 => "000000000000000000000000",
3387 => "000000000000000000000000",
3388 => "000000000000000000000000",
3389 => "000000000000000000000000",
3390 => "000000000000000000000000",
3391 => "000000000000000000000000",
3392 => "000000000000000000000000",
3393 => "000000000000000000000000",
3394 => "000000000000000000000000",
3395 => "000000000000000000000000",
3396 => "000000000000000000000000",
3397 => "000000000000000000000000",
3398 => "000000000000000000000000",
3399 => "000000000000000000000000",
3400 => "001101000011010000110100",
3401 => "010100110101001101010011",
3402 => "010100110101001101010011",
3403 => "010100110101001101010011",
3404 => "010100110101001101010011",
3405 => "000111110001111100011111",
3406 => "000000000000000000000000",
3407 => "000000000000000000000000",
3408 => "000000000000000000000000",
3409 => "000000000000000000000000",
3410 => "000000000000000000000000",
3411 => "000000000000000000000000",
3412 => "000000000000000000000000",
3413 => "000000000000000000000000",
3414 => "000000000000000000000000",
3415 => "000000000000000000000000",
3416 => "000000000000000000000000",
3417 => "000000000000000000000000",
3418 => "000000000000000000000000",
3419 => "000000000000000000000000",
3420 => "000000000000000000000000",
3421 => "000000000000000000000000",
3422 => "000000000000000000000000",
3423 => "000000000000000000000000",
3424 => "000000000000000000000000",
3425 => "000000000000000000000000",
3426 => "000110110001101100011011",
3427 => "010010100100101001001010",
3428 => "010100110101001101010011",
3429 => "001101100011011000110110",
3430 => "000011000000110000001100",
3431 => "000000000000000000000000",
3432 => "000101010001010100010101",
3433 => "101101011011010110110101",
3434 => "000101000001010000010100",
3435 => "101000111010001110100011",
3436 => "001001110010011100100111",
3437 => "000101100001011000010110",
3438 => "011001010110010101100101",
3439 => "011100010111000101110001",
3440 => "000011110000111100001111",
3441 => "000000000000000000000000",
3442 => "000000000000000000000000",
3443 => "000000000000000000000000",
3444 => "000000000000000000000000",
3445 => "000000000000000000000000",
3446 => "000000000000000000000000",
3447 => "000000000000000000000000",
3448 => "000000000000000000000000",
3449 => "000000000000000000000000",
3450 => "000000000000000000000000",
3451 => "000000000000000000000000",
3452 => "000000000000000000000000",
3453 => "000000000000000000000000",
3454 => "000000000000000000000000",
3455 => "000000000000000000000000",
3456 => "000000000000000000000000",
3457 => "000000000000000000000000",
3458 => "000000000000000000000000",
3459 => "000000000000000000000000",
3460 => "000000000000000000000000",
3461 => "000000000000000000000000",
3462 => "000000000000000000000000",
3463 => "000000000000000000000000",
3464 => "000000000000000000000000",
3465 => "000000000000000000000000",
3466 => "000000000000000000000000",
3467 => "000000000000000000000000",
3468 => "000000000000000000000000",
3469 => "000000000000000000000000",
3470 => "000000000000000000000000",
3471 => "000000000000000000000000",
3472 => "000000000000000000000000",
3473 => "000000000000000000000000",
3474 => "000000000000000000000000",
3475 => "000000000000000000000000",
3476 => "000000000000000000000000",
3477 => "000000000000000000000000",
3478 => "000000000000000000000000",
3479 => "000000000000000000000000",
3480 => "000000000000000000000000",
3481 => "000000000000000000000000",
3482 => "000000000000000000000000",
3483 => "000000000000000000000000",
3484 => "000000000000000000000000",
3485 => "000000000000000000000000",
3486 => "000000000000000000000000",
3487 => "000000000000000000000000",
3488 => "000000000000000000000000",
3489 => "000000000000000000000000",
3490 => "000000000000000000000000",
3491 => "000000000000000000000000",
3492 => "000000000000000000000000",
3493 => "000000000000000000000000",
3494 => "000000000000000000000000",
3495 => "000000000000000000000000",
3496 => "000000000000000000000000",
3497 => "000000000000000000000000",
3498 => "000000000000000000000000",
3499 => "000000000000000000000000",
3500 => "011110000111100001111000",
3501 => "111111111111111111111111",
3502 => "111101001111010011110100",
3503 => "110100111101001111010011",
3504 => "111110101111101011111010",
3505 => "011000000110000001100000",
3506 => "000000000000000000000000",
3507 => "000000110000001100000011",
3508 => "000000100000001000000010",
3509 => "000000000000000000000000",
3510 => "000000000000000000000000",
3511 => "000000000000000000000000",
3512 => "000000000000000000000000",
3513 => "000000000000000000000000",
3514 => "000000000000000000000000",
3515 => "000000000000000000000000",
3516 => "000000000000000000000000",
3517 => "000000000000000000000000",
3518 => "000000000000000000000000",
3519 => "000000000000000000000000",
3520 => "000000000000000000000000",
3521 => "000000000000000000000000",
3522 => "000000000000000000000000",
3523 => "000000000000000000000000",
3524 => "000000000000000000000000",
3525 => "010010100100101001001010",
3526 => "111011111110111111101111",
3527 => "111001101110011011100110",
3528 => "110111001101110011011100",
3529 => "111110101111101011111010",
3530 => "100011101000111010001110",
3531 => "000000000000000000000000",
3532 => "000011110000111100001111",
3533 => "101000111010001110100011",
3534 => "000100100001001000010010",
3535 => "100001111000011110000111",
3536 => "001011100010111000101110",
3537 => "001011010010110100101101",
3538 => "111010011110100111101001",
3539 => "111100011111000111110001",
3540 => "001000000010000000100000",
3541 => "000000000000000000000000",
3542 => "000000000000000000000000",
3543 => "000000000000000000000000",
3544 => "000000000000000000000000",
3545 => "000000000000000000000000",
3546 => "000000000000000000000000",
3547 => "000000000000000000000000",
3548 => "000001100000011000000110",
3549 => "000000000000000000000000",
3550 => "000000000000000000000000",
3551 => "000000000000000000000000",
3552 => "000000000000000000000000",
3553 => "000000000000000000000000",
3554 => "000000000000000000000000",
3555 => "000000000000000000000000",
3556 => "000000000000000000000000",
3557 => "000000000000000000000000",
3558 => "000000000000000000000000",
3559 => "000000000000000000000000",
3560 => "000000000000000000000000",
3561 => "000000000000000000000000",
3562 => "000000000000000000000000",
3563 => "000000000000000000000000",
3564 => "000000000000000000000000",
3565 => "000000000000000000000000",
3566 => "000000000000000000000000",
3567 => "000000000000000000000000",
3568 => "000000000000000000000000",
3569 => "000000000000000000000000",
3570 => "000000000000000000000000",
3571 => "000000000000000000000000",
3572 => "000000000000000000000000",
3573 => "000000000000000000000000",
3574 => "000000000000000000000000",
3575 => "000000000000000000000000",
3576 => "000000000000000000000000",
3577 => "000000000000000000000000",
3578 => "000000000000000000000000",
3579 => "000000000000000000000000",
3580 => "000000000000000000000000",
3581 => "000000000000000000000000",
3582 => "000000000000000000000000",
3583 => "000000000000000000000000",
3584 => "000000000000000000000000",
3585 => "000000000000000000000000",
3586 => "000000000000000000000000",
3587 => "000000000000000000000000",
3588 => "000000000000000000000000",
3589 => "000000000000000000000000",
3590 => "000000000000000000000000",
3591 => "000000000000000000000000",
3592 => "000000000000000000000000",
3593 => "000000000000000000000000",
3594 => "000000000000000000000000",
3595 => "000000000000000000000000",
3596 => "000000000000000000000000",
3597 => "000000000000000000000000",
3598 => "000000000000000000000000",
3599 => "000000000000000000000000",
3600 => "000010010000100100001001",
3601 => "111111111111111111111111",
3602 => "110001001100010011000100",
3603 => "000011010000110100001101",
3604 => "100010011000100110001001",
3605 => "010001100100011001000110",
3606 => "110100001101000011010000",
3607 => "111101011111010111110101",
3608 => "100011011000110110001101",
3609 => "111011011110110111101101",
3610 => "000100110001001100010011",
3611 => "011000100110001001100010",
3612 => "111001101110011011100110",
3613 => "111000001110000011100000",
3614 => "010101000101010001010100",
3615 => "000101010001010100010101",
3616 => "011011010110110101101101",
3617 => "100000011000000110000001",
3618 => "100111111001111110011111",
3619 => "111011111110111111101111",
3620 => "010111110101111101011111",
3621 => "000000000000000000000000",
3622 => "000000000000000000000000",
3623 => "000000000000000000000000",
3624 => "000100010001000100010001",
3625 => "111001101110011011100110",
3626 => "111000101110001011100010",
3627 => "000110010001100100011001",
3628 => "000100000001000000010000",
3629 => "111110001111100011111000",
3630 => "100101011001010110010101",
3631 => "010011110100111101001111",
3632 => "111101011111010111110101",
3633 => "111101001111010011110100",
3634 => "011111110111111101111111",
3635 => "111101101111011011110110",
3636 => "110111011101110111011101",
3637 => "000000000000000000000000",
3638 => "101111111011111110111111",
3639 => "111100011111000111110001",
3640 => "001000000010000000100000",
3641 => "000111010001110100011101",
3642 => "101111001011110010111100",
3643 => "111100011111000111110001",
3644 => "101000011010000110100001",
3645 => "000010010000100100001001",
3646 => "110001111100011111000111",
3647 => "111101011111010111110101",
3648 => "100110101001101010011010",
3649 => "111010101110101011101010",
3650 => "001101110011011100110111",
3651 => "000000000000000000000000",
3652 => "000000000000000000000000",
3653 => "000000000000000000000000",
3654 => "000000000000000000000000",
3655 => "000000000000000000000000",
3656 => "000000000000000000000000",
3657 => "000000000000000000000000",
3658 => "000000000000000000000000",
3659 => "000000000000000000000000",
3660 => "000000000000000000000000",
3661 => "000000000000000000000000",
3662 => "000000000000000000000000",
3663 => "000000000000000000000000",
3664 => "000000000000000000000000",
3665 => "000000000000000000000000",
3666 => "000000000000000000000000",
3667 => "000000000000000000000000",
3668 => "000000000000000000000000",
3669 => "000000000000000000000000",
3670 => "000000000000000000000000",
3671 => "000000000000000000000000",
3672 => "000000000000000000000000",
3673 => "000000000000000000000000",
3674 => "000000000000000000000000",
3675 => "000000000000000000000000",
3676 => "000000000000000000000000",
3677 => "000000000000000000000000",
3678 => "000000000000000000000000",
3679 => "000000000000000000000000",
3680 => "000000000000000000000000",
3681 => "000000000000000000000000",
3682 => "000000000000000000000000",
3683 => "000000000000000000000000",
3684 => "000000000000000000000000",
3685 => "000000000000000000000000",
3686 => "000000000000000000000000",
3687 => "000000000000000000000000",
3688 => "000000000000000000000000",
3689 => "000000000000000000000000",
3690 => "000000000000000000000000",
3691 => "000000000000000000000000",
3692 => "000000000000000000000000",
3693 => "000000000000000000000000",
3694 => "000000000000000000000000",
3695 => "000000000000000000000000",
3696 => "000000000000000000000000",
3697 => "000000000000000000000000",
3698 => "000000000000000000000000",
3699 => "000000000000000000000000",
3700 => "000001110000011100000111",
3701 => "111111111111111111111111",
3702 => "111111011111110111111101",
3703 => "111110001111100011111000",
3704 => "101011001010110010101100",
3705 => "000001100000011000000110",
3706 => "101001011010010110100101",
3707 => "111111111111111111111111",
3708 => "110101011101010111010101",
3709 => "111101111111011111110111",
3710 => "001111100011111000111110",
3711 => "111101111111011111110111",
3712 => "100010101000101010001010",
3713 => "100101001001010010010100",
3714 => "111010111110101111101011",
3715 => "001000100010001000100010",
3716 => "111001001110010011100100",
3717 => "111111001111110011111100",
3718 => "100101001001010010010100",
3719 => "111101011111010111110101",
3720 => "110111011101110111011101",
3721 => "000000000000000000000000",
3722 => "000000000000000000000000",
3723 => "000000000000000000000000",
3724 => "001011000010110000101100",
3725 => "111101101111011011110110",
3726 => "101100111011001110110011",
3727 => "000000000000000000000000",
3728 => "010011110100111101001111",
3729 => "011011000110110001101100",
3730 => "011010010110100101101001",
3731 => "000100000001000000010000",
3732 => "101111011011110110111101",
3733 => "111110111111101111111011",
3734 => "001001110010011100100111",
3735 => "111010001110100011101000",
3736 => "111001001110010011100100",
3737 => "000000000000000000000000",
3738 => "101111111011111110111111",
3739 => "111100011111000111110001",
3740 => "001000100010001000100010",
3741 => "101100111011001110110011",
3742 => "111000101110001011100010",
3743 => "010001010100010101000101",
3744 => "111101111111011111110111",
3745 => "010111100101111001011110",
3746 => "100110101001101010011010",
3747 => "111111111111111111111111",
3748 => "110110001101100011011000",
3749 => "111100001111000011110000",
3750 => "001110010011100100111001",
3751 => "000000000000000000000000",
3752 => "000000000000000000000000",
3753 => "000000000000000000000000",
3754 => "000000000000000000000000",
3755 => "000000000000000000000000",
3756 => "000000000000000000000000",
3757 => "000000000000000000000000",
3758 => "000000000000000000000000",
3759 => "000000000000000000000000",
3760 => "000000000000000000000000",
3761 => "000000000000000000000000",
3762 => "000000000000000000000000",
3763 => "000000000000000000000000",
3764 => "000000000000000000000000",
3765 => "000000000000000000000000",
3766 => "000000000000000000000000",
3767 => "000000000000000000000000",
3768 => "000000000000000000000000",
3769 => "000000000000000000000000",
3770 => "000000000000000000000000",
3771 => "000000000000000000000000",
3772 => "000000000000000000000000",
3773 => "000000000000000000000000",
3774 => "000000000000000000000000",
3775 => "000000000000000000000000",
3776 => "000000000000000000000000",
3777 => "000000000000000000000000",
3778 => "000000000000000000000000",
3779 => "000000000000000000000000",
3780 => "000000000000000000000000",
3781 => "000000000000000000000000",
3782 => "000000000000000000000000",
3783 => "000000000000000000000000",
3784 => "000000000000000000000000",
3785 => "000000000000000000000000",
3786 => "000000000000000000000000",
3787 => "000000000000000000000000",
3788 => "000000000000000000000000",
3789 => "000000000000000000000000",
3790 => "000000000000000000000000",
3791 => "000000000000000000000000",
3792 => "000000000000000000000000",
3793 => "000000000000000000000000",
3794 => "000000000000000000000000",
3795 => "000000000000000000000000",
3796 => "000000000000000000000000",
3797 => "000000000000000000000000",
3798 => "000000000000000000000000",
3799 => "000000000000000000000000",
3800 => "000001110000011100000111",
3801 => "111111111111111111111111",
3802 => "110111011101110111011101",
3803 => "011011000110110001101100",
3804 => "010010110100101101001011",
3805 => "000000000000000000000000",
3806 => "010110000101100001011000",
3807 => "111111111111111111111111",
3808 => "010100010101000101010001",
3809 => "000001000000010000000100",
3810 => "010100100101001001010010",
3811 => "111111111111111111111111",
3812 => "111010001110100011101000",
3813 => "110111111101111111011111",
3814 => "111000011110000111100001",
3815 => "000111010001110100011101",
3816 => "101110101011101010111010",
3817 => "111101111111011111110111",
3818 => "001001010010010100100101",
3819 => "111001101110011011100110",
3820 => "110111111101111111011111",
3821 => "000000000000000000000000",
3822 => "000000000000000000000000",
3823 => "000000000000000000000000",
3824 => "001010010010100100101001",
3825 => "111101011111010111110101",
3826 => "110000011100000111000001",
3827 => "000000110000001100000011",
3828 => "100101111001011110010111",
3829 => "111111101111111011111110",
3830 => "110111011101110111011101",
3831 => "000110010001100100011001",
3832 => "101101111011011110110111",
3833 => "111110111111101111111011",
3834 => "001001000010010000100100",
3835 => "111000111110001111100011",
3836 => "111001001110010011100100",
3837 => "000000000000000000000000",
3838 => "101111111011111110111111",
3839 => "111100011111000111110001",
3840 => "001011010010110100101101",
3841 => "111000111110001111100011",
3842 => "111110001111100011111000",
3843 => "110111101101111011011110",
3844 => "111000011110000111100001",
3845 => "100011011000110110001101",
3846 => "010010010100100101001001",
3847 => "111111101111111011111110",
3848 => "011100000111000001110000",
3849 => "000001000000010000000100",
3850 => "000000010000000100000001",
3851 => "000000000000000000000000",
3852 => "000000000000000000000000",
3853 => "000000000000000000000000",
3854 => "000000000000000000000000",
3855 => "000000000000000000000000",
3856 => "000000000000000000000000",
3857 => "000000000000000000000000",
3858 => "000000000000000000000000",
3859 => "000000000000000000000000",
3860 => "000000000000000000000000",
3861 => "000000000000000000000000",
3862 => "000000000000000000000000",
3863 => "000000000000000000000000",
3864 => "000000000000000000000000",
3865 => "000000000000000000000000",
3866 => "000000000000000000000000",
3867 => "000000000000000000000000",
3868 => "000000000000000000000000",
3869 => "000000000000000000000000",
3870 => "000000000000000000000000",
3871 => "000000000000000000000000",
3872 => "000000000000000000000000",
3873 => "000000000000000000000000",
3874 => "000000000000000000000000",
3875 => "000000000000000000000000",
3876 => "000000000000000000000000",
3877 => "000000000000000000000000",
3878 => "000000000000000000000000",
3879 => "000000000000000000000000",
3880 => "000000000000000000000000",
3881 => "000000000000000000000000",
3882 => "000000000000000000000000",
3883 => "000000000000000000000000",
3884 => "000000000000000000000000",
3885 => "000000000000000000000000",
3886 => "000000000000000000000000",
3887 => "000000000000000000000000",
3888 => "000000000000000000000000",
3889 => "000000000000000000000000",
3890 => "000000000000000000000000",
3891 => "000000000000000000000000",
3892 => "000000000000000000000000",
3893 => "000000000000000000000000",
3894 => "000000000000000000000000",
3895 => "000000000000000000000000",
3896 => "000000000000000000000000",
3897 => "000000000000000000000000",
3898 => "000000000000000000000000",
3899 => "000000000000000000000000",
3900 => "000110000001100000011000",
3901 => "111111111111111111111111",
3902 => "110100001101000011010000",
3903 => "001110110011101100111011",
3904 => "110101101101011011010110",
3905 => "100000011000000110000001",
3906 => "010110000101100001011000",
3907 => "111111111111111111111111",
3908 => "010010100100101001001010",
3909 => "000000000000000000000000",
3910 => "001110000011100000111000",
3911 => "111110111111101111111011",
3912 => "110000001100000011000000",
3913 => "010101000101010001010100",
3914 => "101010001010100010101000",
3915 => "000000010000000100000001",
3916 => "101110101011101010111010",
3917 => "111101111111011111110111",
3918 => "001001010010010100100101",
3919 => "111001101110011011100110",
3920 => "111000011110000111100001",
3921 => "000001000000010000000100",
3922 => "000000000000000000000000",
3923 => "000000000000000000000000",
3924 => "000010100000101000001010",
3925 => "110100101101001011010010",
3926 => "111111001111110011111100",
3927 => "100000101000001010000010",
3928 => "011101010111010101110101",
3929 => "111111011111110111111101",
3930 => "100101011001010110010101",
3931 => "000000000000000000000000",
3932 => "101101111011011110110111",
3933 => "111111011111110111111101",
3934 => "011101110111011101110111",
3935 => "111101111111011111110111",
3936 => "111001001110010011100100",
3937 => "000000000000000000000000",
3938 => "101111111011111110111111",
3939 => "111100011111000111110001",
3940 => "001001000010010000100100",
3941 => "110010111100101111001011",
3942 => "111100011111000111110001",
3943 => "011001110110011101100111",
3944 => "011011100110111001101110",
3945 => "011010000110100001101000",
3946 => "010010010100100101001001",
3947 => "111111101111111011111110",
3948 => "011010010110100101101001",
3949 => "000000000000000000000000",
3950 => "000000000000000000000000",
3951 => "000000000000000000000000",
3952 => "000000000000000000000000",
3953 => "000000000000000000000000",
3954 => "000000000000000000000000",
3955 => "000000000000000000000000",
3956 => "000000000000000000000000",
3957 => "000000000000000000000000",
3958 => "000000000000000000000000",
3959 => "000000000000000000000000",
3960 => "000000000000000000000000",
3961 => "000000000000000000000000",
3962 => "000000000000000000000000",
3963 => "000000000000000000000000",
3964 => "000000000000000000000000",
3965 => "000000000000000000000000",
3966 => "000000000000000000000000",
3967 => "000000000000000000000000",
3968 => "000000000000000000000000",
3969 => "000000000000000000000000",
3970 => "000000000000000000000000",
3971 => "000000000000000000000000",
3972 => "000000000000000000000000",
3973 => "000000000000000000000000",
3974 => "000000000000000000000000",
3975 => "000000000000000000000000",
3976 => "000000000000000000000000",
3977 => "000000000000000000000000",
3978 => "000000000000000000000000",
3979 => "000000000000000000000000",
3980 => "000000000000000000000000",
3981 => "000000000000000000000000",
3982 => "000000000000000000000000",
3983 => "000000000000000000000000",
3984 => "000000000000000000000000",
3985 => "000000000000000000000000",
3986 => "000000000000000000000000",
3987 => "000000000000000000000000",
3988 => "000000000000000000000000",
3989 => "000000000000000000000000",
3990 => "000000000000000000000000",
3991 => "000000000000000000000000",
3992 => "000000000000000000000000",
3993 => "000000000000000000000000",
3994 => "000000000000000000000000",
3995 => "000000000000000000000000",
3996 => "000000000000000000000000",
3997 => "000000000000000000000000",
3998 => "000000000000000000000000",
3999 => "000000000000000000000000",
4000 => "101000001010000010100000",
4001 => "111111111111111111111111",
4002 => "111111111111111111111111",
4003 => "111111101111111011111110",
4004 => "111111111111111111111111",
4005 => "100011001000110010001100",
4006 => "110110001101100011011000",
4007 => "111111111111111111111111",
4008 => "110110101101101011011010",
4009 => "000011000000110000001100",
4010 => "000000110000001100000011",
4011 => "100011111000111110001111",
4012 => "111101001111010011110100",
4013 => "111101011111010111110101",
4014 => "100110001001100010011000",
4015 => "001101110011011100110111",
4016 => "111111111111111111111111",
4017 => "111111111111111111111111",
4018 => "100101001001010010010100",
4019 => "111001101110011011100110",
4020 => "111111111111111111111111",
4021 => "011001100110011001100110",
4022 => "000000000000000000000000",
4023 => "000000000000000000000000",
4024 => "000000000000000000000000",
4025 => "001001000010010000100100",
4026 => "101101101011011010110110",
4027 => "111101111111011111110111",
4028 => "111111111111111111111111",
4029 => "110101101101011011010110",
4030 => "010111010101110101011101",
4031 => "000000000000000000000000",
4032 => "010111110101111101011111",
4033 => "111101111111011111110111",
4034 => "110010101100101011001010",
4035 => "111010001110100011101000",
4036 => "111111111111111111111111",
4037 => "011011010110110101101101",
4038 => "111111111111111111111111",
4039 => "111111111111111111111111",
4040 => "100110111001101110011011",
4041 => "001101010011010100110101",
4042 => "110110001101100011011000",
4043 => "111111101111111011111110",
4044 => "110010001100100011001000",
4045 => "001101100011011000110110",
4046 => "110011111100111111001111",
4047 => "111111111111111111111111",
4048 => "111111101111111011111110",
4049 => "000000000000000000000000",
4050 => "000000000000000000000000",
4051 => "000000000000000000000000",
4052 => "000000000000000000000000",
4053 => "000000000000000000000000",
4054 => "000000000000000000000000",
4055 => "000000000000000000000000",
4056 => "000000000000000000000000",
4057 => "000000000000000000000000",
4058 => "000000000000000000000000",
4059 => "000000000000000000000000",
4060 => "000000000000000000000000",
4061 => "000000000000000000000000",
4062 => "000000000000000000000000",
4063 => "000000000000000000000000",
4064 => "000000000000000000000000",
4065 => "000000000000000000000000",
4066 => "000000000000000000000000",
4067 => "000000000000000000000000",
4068 => "000000000000000000000000",
4069 => "000000000000000000000000",
4070 => "000000000000000000000000",
4071 => "000000000000000000000000",
4072 => "000000000000000000000000",
4073 => "000000000000000000000000",
4074 => "000000000000000000000000",
4075 => "000000000000000000000000",
4076 => "000000000000000000000000",
4077 => "000000000000000000000000",
4078 => "000000000000000000000000",
4079 => "000000000000000000000000",
4080 => "000000000000000000000000",
4081 => "000000000000000000000000",
4082 => "000000000000000000000000",
4083 => "000000000000000000000000",
4084 => "000000000000000000000000",
4085 => "000000000000000000000000",
4086 => "000000000000000000000000",
4087 => "000000000000000000000000",
4088 => "000000000000000000000000",
4089 => "000000000000000000000000",
4090 => "000000000000000000000000",
4091 => "000000000000000000000000",
4092 => "000000000000000000000000",
4093 => "000000000000000000000000",
4094 => "000000000000000000000000",
4095 => "000000000000000000000000",
4096 => "000000000000000000000000",
4097 => "000000000000000000000000",
4098 => "000000000000000000000000",
4099 => "000000000000000000000000",
4100 => "000000000000000000000000",
4101 => "000000000000000000000000",
4102 => "000000000000000000000000",
4103 => "000000000000000000000000",
4104 => "000000000000000000000000",
4105 => "000000000000000000000000",
4106 => "000000000000000000000000",
4107 => "000000000000000000000000",
4108 => "000000000000000000000000",
4109 => "000000000000000000000000",
4110 => "000000000000000000000000",
4111 => "000000000000000000000000",
4112 => "000000000000000000000000",
4113 => "000000000000000000000000",
4114 => "000000000000000000000000",
4115 => "000000000000000000000000",
4116 => "000000000000000000000000",
4117 => "000000000000000000000000",
4118 => "000000000000000000000000",
4119 => "000000000000000000000000",
4120 => "000000000000000000000000",
4121 => "000000000000000000000000",
4122 => "000000000000000000000000",
4123 => "000000000000000000000000",
4124 => "000000000000000000000000",
4125 => "000000000000000000000000",
4126 => "000000000000000000000000",
4127 => "000000000000000000000000",
4128 => "000000000000000000000000",
4129 => "000000000000000000000000",
4130 => "000000000000000000000000",
4131 => "000000000000000000000000",
4132 => "000000000000000000000000",
4133 => "000000000000000000000000",
4134 => "000000010000000100000001",
4135 => "000110010001100100011001",
4136 => "000010010000100100001001",
4137 => "000000000000000000000000",
4138 => "000000000000000000000000",
4139 => "000000000000000000000000",
4140 => "000000000000000000000000",
4141 => "000000000000000000000000",
4142 => "000000000000000000000000",
4143 => "000000000000000000000000",
4144 => "000000000000000000000000",
4145 => "000000000000000000000000",
4146 => "000000000000000000000000",
4147 => "000000000000000000000000",
4148 => "000000000000000000000000",
4149 => "000000000000000000000000",
4150 => "000000000000000000000000",
4151 => "000000000000000000000000",
4152 => "000000000000000000000000",
4153 => "000000000000000000000000",
4154 => "000000000000000000000000",
4155 => "000000000000000000000000",
4156 => "000000000000000000000000",
4157 => "000000000000000000000000",
4158 => "000000000000000000000000",
4159 => "000000000000000000000000",
4160 => "000000000000000000000000",
4161 => "000000000000000000000000",
4162 => "000000000000000000000000",
4163 => "000000000000000000000000",
4164 => "000000000000000000000000",
4165 => "000000000000000000000000",
4166 => "000000000000000000000000",
4167 => "000000000000000000000000",
4168 => "000000000000000000000000",
4169 => "000000000000000000000000",
4170 => "000000000000000000000000",
4171 => "000000000000000000000000",
4172 => "000000000000000000000000",
4173 => "000000000000000000000000",
4174 => "000000000000000000000000",
4175 => "000000000000000000000000",
4176 => "000000000000000000000000",
4177 => "000000000000000000000000",
4178 => "000000000000000000000000",
4179 => "000000000000000000000000",
4180 => "000000000000000000000000",
4181 => "000000000000000000000000",
4182 => "000000000000000000000000",
4183 => "000000000000000000000000",
4184 => "000000000000000000000000",
4185 => "000000000000000000000000",
4186 => "000000000000000000000000",
4187 => "000000000000000000000000",
4188 => "000000000000000000000000",
4189 => "000000000000000000000000",
4190 => "000000000000000000000000",
4191 => "000000000000000000000000",
4192 => "000000000000000000000000",
4193 => "000000000000000000000000",
4194 => "000000000000000000000000",
4195 => "000000000000000000000000",
4196 => "000000000000000000000000",
4197 => "000000000000000000000000",
4198 => "000000000000000000000000",
4199 => "000000000000000000000000"

    );
begin
    data_out <= ROM_Data(to_integer(unsigned(address)));
end architecture Behavioral;