library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;
use ieee.numeric_std.all;

entity alienship is
    Port (
        address : in STD_LOGIC_VECTOR(13 downto 0);
        data_out : out STD_LOGIC_VECTOR(23 downto 0)
    );
end entity alienship;

architecture Behavioral of alienship is
    type ROM_Type is array (0 to 4899) of STD_LOGIC_VECTOR(23 downto 0);
    constant ROM_Data : ROM_Type := (
0 => "000000000000000000000000",
1 => "000000000000000000000000",
2 => "000000000000000000000000",
3 => "000000000000000000000000",
4 => "000000000000000000000000",
5 => "000000000000000000000000",
6 => "000000000000000000000000",
7 => "000000000000000000000000",
8 => "000000000000000000000000",
9 => "000000000000000000000000",
10 => "000000000000000000000000",
11 => "000000000000000000000000",
12 => "000000000000000000000000",
13 => "000000000000000000000000",
14 => "000000000000000000000000",
15 => "000000000000000000000000",
16 => "000000000000000000000000",
17 => "000000000000000000000000",
18 => "000000000000000000000000",
19 => "000000000000000000000000",
20 => "000000110000000100000010",
21 => "000001010000001100000100",
22 => "000000000000000000000000",
23 => "000000000000000000000000",
24 => "000000000000000000000000",
25 => "000000000000000000000000",
26 => "000000000000000000000000",
27 => "000000000000000000000000",
28 => "000000000000000000000000",
29 => "000000000000000000000000",
30 => "000000000000000000000000",
31 => "000000000000000000000000",
32 => "000000000000000000000000",
33 => "000000000000000000000000",
34 => "000000000000000000000000",
35 => "000000000000000000000000",
36 => "000000000000000000000000",
37 => "000001000000001000011000",
38 => "000000010000000000000110",
39 => "000000000000000000000000",
40 => "000000000000000000000000",
41 => "000000000000000000000000",
42 => "000000000000000000000000",
43 => "000000000000000000000000",
44 => "000000000000000000000000",
45 => "000000000000000000000000",
46 => "000000000000000000000000",
47 => "000000000000000000000000",
48 => "000000000000000000000000",
49 => "000000000000000000000000",
50 => "000000000000000000000000",
51 => "000000000000000000000000",
52 => "000000000000000000000000",
53 => "000000000000000000000000",
54 => "000001000000001000000011",
55 => "000000110000001000000010",
56 => "000000000000000000000000",
57 => "000000000000000000000000",
58 => "000000000000000000000000",
59 => "000000000000000000000000",
60 => "000000000000000000000000",
61 => "000000000000000000000000",
62 => "000000000000000000000000",
63 => "000000000000000000000000",
64 => "000000000000000000000000",
65 => "000000000000000000000000",
66 => "000000000000000000000000",
67 => "000000000000000000000000",
68 => "000000000000000000000000",
69 => "000000000000000000000000",
70 => "000000000000000000000000",
71 => "000000000000000000000000",
72 => "000000000000000000000000",
73 => "000000000000000000000000",
74 => "000000000000000000000000",
75 => "000000000000000000000000",
76 => "000000000000000000000000",
77 => "000000000000000000000000",
78 => "000000000000000000000000",
79 => "000000000000000000000000",
80 => "000000000000000000000000",
81 => "000000000000000000000000",
82 => "000000000000000000000000",
83 => "000000000000000000000000",
84 => "000000000000000000000000",
85 => "000000000000000000000000",
86 => "000000000000000000000000",
87 => "000000000000000000000000",
88 => "000000000000000000000000",
89 => "000000000000000000000000",
90 => "000111110010001100100100",
91 => "000011000000101100001100",
92 => "000000000000000000000000",
93 => "000000000000000000000000",
94 => "000000000000000000000000",
95 => "000000000000000000000000",
96 => "000000000000000000000000",
97 => "000000000000000000000000",
98 => "000000000000000000000000",
99 => "000000000000000000000000",
100 => "000000000000000000000000",
101 => "000000000000000000000000",
102 => "000000000000000000000000",
103 => "000000000000000000000000",
104 => "000000000000000000000000",
105 => "000000000000000000000000",
106 => "000000000000000000000000",
107 => "000000110000000100011011",
108 => "000001010000001100100000",
109 => "000000000000000000000000",
110 => "000000000000000000000000",
111 => "000000000000000000000000",
112 => "000000000000000000000000",
113 => "000000000000000000000000",
114 => "000000000000000000000000",
115 => "000000000000000000000000",
116 => "000000000000000000000000",
117 => "000000000000000000000000",
118 => "000000000000000000000000",
119 => "000000000000000000000000",
120 => "000000000000000000000000",
121 => "000000000000000000000000",
122 => "000000000000000000000000",
123 => "000000000000000000000000",
124 => "000010110000101000001011",
125 => "001001000010010100100111",
126 => "000000010000000100000001",
127 => "000000000000000000000000",
128 => "000000000000000000000000",
129 => "000000000000000000000000",
130 => "000000000000000000000000",
131 => "000000000000000000000000",
132 => "000000000000000000000000",
133 => "000000000000000000000000",
134 => "000000000000000000000000",
135 => "000000000000000000000000",
136 => "000000000000000000000000",
137 => "000000000000000000000000",
138 => "000000000000000000000000",
139 => "000000000000000000000000",
140 => "000000000000000000000000",
141 => "000000000000000000000000",
142 => "000000000000000000000000",
143 => "000000000000000000000000",
144 => "000000000000000000000000",
145 => "000000000000000000000000",
146 => "000000000000000000000000",
147 => "000000000000000000000000",
148 => "000000000000000000000000",
149 => "000000000000000000000000",
150 => "000000000000000000000000",
151 => "000000000000000000000000",
152 => "000000000000000000000000",
153 => "000000000000000000000000",
154 => "000000000000000000000000",
155 => "000000000000000000000000",
156 => "000000000000000000000000",
157 => "000000000000000000000000",
158 => "000000000000000000000000",
159 => "000001110000011000000111",
160 => "001000000010010100100101",
161 => "000000000000000000000000",
162 => "000000000000000000000000",
163 => "000000000000000000000000",
164 => "000000000000000000000000",
165 => "000000000000000000000000",
166 => "000000000000000000000000",
167 => "000000000000000000000000",
168 => "000000000000000000000000",
169 => "000000000000000000000000",
170 => "000000000000000000000000",
171 => "000000000000000000000000",
172 => "000000000000000000000000",
173 => "000000000000000000000000",
174 => "000000000000000000000000",
175 => "000000000000000000000000",
176 => "000000000000000000000000",
177 => "000001010000001000100100",
178 => "000000100000001000011001",
179 => "000000000000000000000000",
180 => "000000000000000000000000",
181 => "000000000000000000000000",
182 => "000000000000000000000000",
183 => "000000000000000000000000",
184 => "000000000000000000000000",
185 => "000000000000000000000000",
186 => "000000000000000000000000",
187 => "000000000000000000000000",
188 => "000000000000000000000000",
189 => "000000000000000000000000",
190 => "000000000000000000000000",
191 => "000000000000000000000000",
192 => "000000000000000000000000",
193 => "000000000000000000000000",
194 => "000000000000000000000000",
195 => "000111100010010100100101",
196 => "000001110000100000001001",
197 => "000000000000000000000000",
198 => "000000000000000000000000",
199 => "000000000000000000000000",
200 => "000000000000000000000000",
201 => "000000000000000000000000",
202 => "000000000000000000000000",
203 => "000000000000000000000000",
204 => "000000000000000000000000",
205 => "000000000000000000000000",
206 => "000000000000000000000000",
207 => "000000000000000000000000",
208 => "000000000000000000000000",
209 => "000000000000000000000000",
210 => "000000000000000000000000",
211 => "000000000000000000000000",
212 => "000000000000000000000000",
213 => "000000000000000000000000",
214 => "000000000000000000000000",
215 => "000000000000000000000000",
216 => "000000000000000000000000",
217 => "000000000000000000000000",
218 => "000000000000000000000000",
219 => "000000000000000000000000",
220 => "000000000000000000000000",
221 => "000000000000000000000000",
222 => "000000000000000000000000",
223 => "000000000000000000000000",
224 => "000000000000000000000000",
225 => "000000000000000000000000",
226 => "000000000000000000000000",
227 => "000000000000000000000000",
228 => "000000000000000000000000",
229 => "000011010001000000001111",
230 => "000101110001011100010111",
231 => "000000000000000000000000",
232 => "000000000000000000000000",
233 => "000000000000000000000000",
234 => "000000000000000000000000",
235 => "000000000000000000000000",
236 => "000000000000000000000000",
237 => "000000000000000000000000",
238 => "000000000000000000000000",
239 => "000000000000000000000000",
240 => "000000000000000000000000",
241 => "000000000000000000000000",
242 => "000000000000000000000000",
243 => "000000000000000000000000",
244 => "000000000000000000000000",
245 => "000000000000000000000000",
246 => "000000000000000000000000",
247 => "000001100000001000110100",
248 => "000000100000001100100011",
249 => "000000000000000000000000",
250 => "000000000000000000000000",
251 => "000000000000000000000000",
252 => "000000000000000000000000",
253 => "000000000000000000000000",
254 => "000000000000000000000000",
255 => "000000000000000000000000",
256 => "000000000000000000000000",
257 => "000000000000000000000000",
258 => "000000000000000000000000",
259 => "000000000000000000000000",
260 => "000000000000000000000000",
261 => "000000000000000000000000",
262 => "000000000000000000000000",
263 => "000000000000000000000000",
264 => "000000000000000000000000",
265 => "000100100001011000010110",
266 => "000011110001000100010001",
267 => "000000000000000000000000",
268 => "000000000000000000000000",
269 => "000000000000000000000000",
270 => "000000000000000000000000",
271 => "000000000000000000000000",
272 => "000000000000000000000000",
273 => "000000000000000000000000",
274 => "000000000000000000000000",
275 => "000000000000000000000000",
276 => "000000000000000000000000",
277 => "000000000000000000000000",
278 => "000000000000000000000000",
279 => "000000000000000000000000",
280 => "000000000000000000000000",
281 => "000000000000000000000000",
282 => "000000000000000000000000",
283 => "000000000000000000000000",
284 => "000000000000000000000000",
285 => "000000000000000000000000",
286 => "000000000000000000000000",
287 => "000000000000000000000000",
288 => "000000000000000000000000",
289 => "000000000000000000000000",
290 => "000000000000000000000000",
291 => "000000000000000000000000",
292 => "000000000000000000000000",
293 => "000000000000000000000000",
294 => "000000000000000000000000",
295 => "000000000000000000000000",
296 => "000000000000000000000000",
297 => "000000000000000000000000",
298 => "000000000000000000000000",
299 => "000110010001100000011000",
300 => "000001000000001000000011",
301 => "000000000000000000000000",
302 => "000000000000000000000000",
303 => "000000000000000000000000",
304 => "000000000000000000000000",
305 => "000000000000000000000000",
306 => "000000000000000000000000",
307 => "000000000000000000000000",
308 => "000000000000000000000000",
309 => "000000000000000000000000",
310 => "000000000000000000000000",
311 => "000000000000000000000000",
312 => "000000000000000000000000",
313 => "000000000000000000000000",
314 => "000000000000000000000000",
315 => "000000000000000000000000",
316 => "000000000000000000000000",
317 => "000001000000001000110111",
318 => "000000110000001100111100",
319 => "000000000000000000000000",
320 => "000000000000000000000000",
321 => "000000000000000000000000",
322 => "000000000000000000000000",
323 => "000000000000000000000000",
324 => "000000000000000000000000",
325 => "000000000000000000000000",
326 => "000000000000000000000000",
327 => "000000000000000000000000",
328 => "000000000000000000000000",
329 => "000000000000000000000000",
330 => "000000000000000000000000",
331 => "000000000000000000000000",
332 => "000000000000000000000000",
333 => "000000000000000000000000",
334 => "000000000000000000000000",
335 => "000000010000000100000001",
336 => "000111100001101100011011",
337 => "000000000000000000000000",
338 => "000000000000000000000000",
339 => "000000000000000000000000",
340 => "000000000000000000000000",
341 => "000000000000000000000000",
342 => "000000000000000000000000",
343 => "000000000000000000000000",
344 => "000000000000000000000000",
345 => "000000000000000000000000",
346 => "000000000000000000000000",
347 => "000000000000000000000000",
348 => "000000000000000000000000",
349 => "000000000000000000000000",
350 => "000000000000000000000000",
351 => "000000000000000000000000",
352 => "000000000000000000000000",
353 => "000000000000000000000000",
354 => "000000000000000000000000",
355 => "000000000000000000000000",
356 => "000000000000000000000000",
357 => "000000000000000000000000",
358 => "000000000000000000000000",
359 => "000000000000000000000000",
360 => "000000000000000000000000",
361 => "000000000000000000000000",
362 => "000000000000000000000000",
363 => "000000000000000000000000",
364 => "000000000000000000000000",
365 => "000000000000000000000000",
366 => "000000000000000000000000",
367 => "000000000000000000000000",
368 => "000000100000000100000010",
369 => "000101100001001000010010",
370 => "000000100000000100000001",
371 => "000000000000000000000000",
372 => "000000000000000000000000",
373 => "000000000000000000000000",
374 => "000000000000000000000000",
375 => "000000000000000000000000",
376 => "000000000000000000000000",
377 => "000000000000000000000000",
378 => "000000000000000000000000",
379 => "000000000000000000000000",
380 => "000000000000000000000000",
381 => "000000000000000000000000",
382 => "000000000000000000000000",
383 => "000000000000000000000000",
384 => "000000000000000000000000",
385 => "000000000000000000000001",
386 => "000001010000010000010111",
387 => "000001000000001100111111",
388 => "000001000000001100111111",
389 => "000001100000010000011111",
390 => "000000000000000000000000",
391 => "000000000000000000000000",
392 => "000000000000000000000000",
393 => "000000000000000000000000",
394 => "000000000000000000000000",
395 => "000000000000000000000000",
396 => "000000000000000000000000",
397 => "000000000000000000000000",
398 => "000000000000000000000000",
399 => "000000000000000000000000",
400 => "000000000000000000000000",
401 => "000000000000000000000000",
402 => "000000000000000000000000",
403 => "000000000000000000000000",
404 => "000000000000000000000000",
405 => "000000000000000000000000",
406 => "000100110001000100001111",
407 => "000000100000001000000010",
408 => "000000000000000000000000",
409 => "000000000000000000000000",
410 => "000000000000000000000000",
411 => "000000000000000000000000",
412 => "000000000000000000000000",
413 => "000000000000000000000000",
414 => "000000000000000000000000",
415 => "000000000000000000000000",
416 => "000000000000000000000000",
417 => "000000000000000000000000",
418 => "000000000000000000000000",
419 => "000000000000000000000000",
420 => "000000000000000000000000",
421 => "000000000000000000000000",
422 => "000000000000000000000000",
423 => "000000000000000000000000",
424 => "000000000000000000000000",
425 => "000000000000000000000000",
426 => "000000000000000000000000",
427 => "000000000000000000000000",
428 => "000000000000000000000000",
429 => "000000000000000000000000",
430 => "000000000000000000000000",
431 => "000000000000000000000000",
432 => "000000000000000000000000",
433 => "000000000000000000000000",
434 => "000000000000000000000000",
435 => "000000000000000000000000",
436 => "000000000000000000000000",
437 => "000000000000000000000000",
438 => "000001010000001000000011",
439 => "000110100001011000010111",
440 => "000000000000000000000000",
441 => "000000000000000000000000",
442 => "000000000000000000000000",
443 => "000000000000000000000000",
444 => "000000000000000000000000",
445 => "000000000000000000000000",
446 => "000000000000000000000000",
447 => "000000000000000000000000",
448 => "000000000000000000000000",
449 => "000000000000000000000000",
450 => "000000000000000000000000",
451 => "000000000000000000000000",
452 => "000000000000000000000000",
453 => "000000000000000000000000",
454 => "000000000000000000000000",
455 => "000000000000000000000100",
456 => "000100010000111010000100",
457 => "000010000000011110011111",
458 => "000001110000101010011110",
459 => "000100000000111110000000",
460 => "000000000000000000000001",
461 => "000000000000000000000000",
462 => "000000000000000000000000",
463 => "000000000000000000000000",
464 => "000000000000000000000000",
465 => "000000000000000000000000",
466 => "000000000000000000000000",
467 => "000000000000000000000000",
468 => "000000000000000000000000",
469 => "000000000000000000000000",
470 => "000000000000000000000000",
471 => "000000000000000000000000",
472 => "000000000000000000000000",
473 => "000000000000000000000000",
474 => "000000000000000000000000",
475 => "000000000000000000000000",
476 => "000101010001010000010010",
477 => "000001010000010000000100",
478 => "000000000000000000000000",
479 => "000000000000000000000000",
480 => "000000000000000000000000",
481 => "000000000000000000000000",
482 => "000000000000000000000000",
483 => "000000000000000000000000",
484 => "000000000000000000000000",
485 => "000000000000000000000000",
486 => "000000000000000000000000",
487 => "000000000000000000000000",
488 => "000000000000000000000000",
489 => "000000000000000000000000",
490 => "000000000000000000000000",
491 => "000000000000000000000000",
492 => "000000000000000000000000",
493 => "000000000000000000000000",
494 => "000000000000000000000000",
495 => "000000000000000000000000",
496 => "000000000000000000000000",
497 => "000000000000000000000000",
498 => "000000000000000000000000",
499 => "000000000000000000000000",
500 => "000000000000000000000000",
501 => "000000000000000000000000",
502 => "000000000000000000000000",
503 => "000000000000000000000000",
504 => "000000000000000000000000",
505 => "000000000000000000000000",
506 => "000000000000000000000000",
507 => "000000000000000000000000",
508 => "000010010000011000000111",
509 => "000100110000111100010001",
510 => "000000000000000000000000",
511 => "000000000000000000000000",
512 => "000000000000000000000000",
513 => "000000000000000000000000",
514 => "000000000000000000000000",
515 => "000000000000000000000000",
516 => "000000000000000000000000",
517 => "000000000000000000000000",
518 => "000000000000000000000000",
519 => "000000000000000000000000",
520 => "000000000000000000000000",
521 => "000000000000000000000000",
522 => "000000000000000000000000",
523 => "000000000000000000000000",
524 => "000000000000000000000000",
525 => "000000000000000000000011",
526 => "000011110001000010001100",
527 => "000010110000110110111110",
528 => "000010010000110010111100",
529 => "000011110001000010001110",
530 => "000000000000000000000010",
531 => "000000000000000000000000",
532 => "000000000000000000000000",
533 => "000000000000000000000000",
534 => "000000000000000000000000",
535 => "000000000000000000000000",
536 => "000000000000000000000000",
537 => "000000000000000000000000",
538 => "000000000000000000000000",
539 => "000000000000000000000000",
540 => "000000000000000000000000",
541 => "000000000000000000000000",
542 => "000000000000000000000000",
543 => "000000000000000000000000",
544 => "000000000000000000000000",
545 => "000000000000000000000000",
546 => "000011100000110100001100",
547 => "000010010000100000000111",
548 => "000000000000000000000000",
549 => "000000000000000000000000",
550 => "000000000000000000000000",
551 => "000000000000000000000000",
552 => "000000000000000000000000",
553 => "000000000000000000000000",
554 => "000000000000000000000000",
555 => "000000000000000000000000",
556 => "000000000000000000000000",
557 => "000000000000000000000000",
558 => "000000000000000000000000",
559 => "000000000000000000000000",
560 => "000000000000000000000000",
561 => "000000000000000000000000",
562 => "000000000000000000000000",
563 => "000000000000000000000000",
564 => "000000000000000000000000",
565 => "000000000000000000000000",
566 => "000000000000000000000000",
567 => "000000000000000000000000",
568 => "000000000000000000000000",
569 => "000000000000000000000000",
570 => "000000000000000000000000",
571 => "000000000000000000000000",
572 => "000000000000000000000000",
573 => "000000000000000000000000",
574 => "000000000000000000000000",
575 => "000000000000000000000000",
576 => "000000000000000000000000",
577 => "000000000000000000000000",
578 => "000100110000111100010000",
579 => "000001110000010000000101",
580 => "000000000000000000000000",
581 => "000000000000000000000000",
582 => "000000000000000000000000",
583 => "000000000000000000000000",
584 => "000000000000000000000000",
585 => "000000000000000000000000",
586 => "000000000000000000000000",
587 => "000000000000000000000000",
588 => "000000000000000000000000",
589 => "000000000000000000000000",
590 => "000000000000000000000000",
591 => "000000000000000000000000",
592 => "000000000000000000000000",
593 => "000000000000000000000000",
594 => "000000000000000000000000",
595 => "000000000000000000000001",
596 => "000010110000101001100011",
597 => "000010110000111010111011",
598 => "000011000000110011000001",
599 => "000011000000101001100001",
600 => "000000000000000000000001",
601 => "000000000000000000000000",
602 => "000000000000000000000000",
603 => "000000000000000000000000",
604 => "000000000000000000000000",
605 => "000000000000000000000000",
606 => "000000000000000000000000",
607 => "000000000000000000000000",
608 => "000000000000000000000000",
609 => "000000000000000000000000",
610 => "000000000000000000000000",
611 => "000000000000000000000000",
612 => "000000000000000000000000",
613 => "000000000000000000000000",
614 => "000000000000000000000000",
615 => "000000000000000000000000",
616 => "000001000000001100000100",
617 => "000101000001000100010001",
618 => "000000000000000000000000",
619 => "000000000000000000000000",
620 => "000000000000000000000000",
621 => "000000000000000000000000",
622 => "000000000000000000000000",
623 => "000000000000000000000000",
624 => "000000000000000000000000",
625 => "000000000000000000000000",
626 => "000000000000000000000000",
627 => "000000000000000000000000",
628 => "000000000000000000000000",
629 => "000000000000000000000000",
630 => "000000000000000000000000",
631 => "000000000000000000000000",
632 => "000000000000000000000000",
633 => "000000000000000000000000",
634 => "000000000000000000000000",
635 => "000000000000000000000000",
636 => "000000000000000000000000",
637 => "000000000000000000000000",
638 => "000000000000000000000000",
639 => "000000000000000000000000",
640 => "000000000000000000000000",
641 => "000000000000000000000000",
642 => "000000000000000000000000",
643 => "000000000000000000000000",
644 => "000000000000000000000000",
645 => "000000000000000000000000",
646 => "000000000000000000000000",
647 => "000000000000000000000000",
648 => "000100010000111000001110",
649 => "000001010000001100000100",
650 => "000000000000000000000000",
651 => "000000000000000000000000",
652 => "000000000000000000000000",
653 => "000000000000000000000000",
654 => "000000000000000000000000",
655 => "000000000000000000000000",
656 => "000000000000000000000000",
657 => "000000000000000000000000",
658 => "000000000000000000000000",
659 => "000000000000000000000000",
660 => "000000000000000000000000",
661 => "000000000000000000000000",
662 => "000000000000000000000000",
663 => "000000000000000000000000",
664 => "000000000000000000000000",
665 => "000001100000010100001011",
666 => "000001000000001100100000",
667 => "000011000000101110011110",
668 => "000011010000101010011100",
669 => "000000110000001100010111",
670 => "000001010000010000001000",
671 => "000000000000000000000000",
672 => "000000000000000000000000",
673 => "000000000000000000000000",
674 => "000000000000000000000000",
675 => "000000000000000000000000",
676 => "000000000000000000000000",
677 => "000000000000000000000000",
678 => "000000000000000000000000",
679 => "000000000000000000000000",
680 => "000000000000000000000000",
681 => "000000000000000000000000",
682 => "000000000000000000000000",
683 => "000000000000000000000000",
684 => "000000000000000000000000",
685 => "000000000000000000000000",
686 => "000000110000001000000011",
687 => "000100110001000000001111",
688 => "000000010000000000000000",
689 => "000000000000000000000000",
690 => "000000000000000000000000",
691 => "000000000000000000000000",
692 => "000000000000000000000000",
693 => "000000000000000000000000",
694 => "000000000000000000000000",
695 => "000000000000000000000000",
696 => "000000000000000000000000",
697 => "000000000000000000000000",
698 => "000000000000000000000000",
699 => "000000000000000000000000",
700 => "000000000000000000000000",
701 => "000000000000000000000000",
702 => "000000000000000000000000",
703 => "000000000000000000000000",
704 => "000000000000000000000000",
705 => "000000000000000000000000",
706 => "000000000000000000000000",
707 => "000000000000000000000000",
708 => "000000000000000000000000",
709 => "000000000000000000000000",
710 => "000000000000000000000000",
711 => "000000000000000000000000",
712 => "000000000000000000000000",
713 => "000000000000000000000000",
714 => "000000000000000000000000",
715 => "000000000000000000000000",
716 => "000000000000000000000000",
717 => "000000100000000100000010",
718 => "000110000001001100010100",
719 => "000000010000000100000001",
720 => "000000000000000000000000",
721 => "000000000000000000000000",
722 => "000000000000000000000000",
723 => "000000000000000000000000",
724 => "000000000000000000000000",
725 => "000000000000000000000000",
726 => "000000000000000000000000",
727 => "000000000000000000000000",
728 => "000000000000000000000000",
729 => "000000000000000000000000",
730 => "000000000000000000000000",
731 => "000000000000000000000000",
732 => "000000000000000000000000",
733 => "000000000000000000000000",
734 => "000000000000000000000000",
735 => "001011100010110001110010",
736 => "000111110010010101100101",
737 => "000100010001001101101000",
738 => "000100010001000101011010",
739 => "001000010010010001011110",
740 => "001011000010110101101101",
741 => "000000000000000000000000",
742 => "000000000000000000000000",
743 => "000000000000000000000000",
744 => "000000000000000000000000",
745 => "000000000000000000000000",
746 => "000000000000000000000000",
747 => "000000000000000000000000",
748 => "000000000000000000000000",
749 => "000000000000000000000000",
750 => "000000000000000000000000",
751 => "000000000000000000000000",
752 => "000000000000000000000000",
753 => "000000000000000000000000",
754 => "000000000000000000000000",
755 => "000000000000000000000000",
756 => "000000010000000100000001",
757 => "000101110001001100010011",
758 => "000000100000001000000010",
759 => "000000000000000000000000",
760 => "000000000000000000000000",
761 => "000000000000000000000000",
762 => "000000000000000000000000",
763 => "000000000000000000000000",
764 => "000000000000000000000000",
765 => "000000000000000000000000",
766 => "000000000000000000000000",
767 => "000000000000000000000000",
768 => "000000000000000000000000",
769 => "000000000000000000000000",
770 => "000000000000000000000000",
771 => "000000000000000000000000",
772 => "000000000000000000000000",
773 => "000000000000000000000000",
774 => "000000000000000000000000",
775 => "000000000000000000000000",
776 => "000000000000000000000000",
777 => "000000000000000000000000",
778 => "000000000000000000000000",
779 => "000000000000000000000000",
780 => "000000000000000000000000",
781 => "000000000000000000000000",
782 => "000000000000000000000000",
783 => "000000000000000000000000",
784 => "000000000000000000000000",
785 => "000000000000000000000000",
786 => "000000000000000000000000",
787 => "000000100000000100000010",
788 => "000110010001010100010101",
789 => "000000000000000000000000",
790 => "000000000000000000000000",
791 => "000000000000000000000000",
792 => "000000000000000000000000",
793 => "000000000000000000000000",
794 => "000000000000000000000000",
795 => "000000000000000000000000",
796 => "000000000000000000000000",
797 => "000000000000000000000000",
798 => "000000000000000000000000",
799 => "000000000000000000000000",
800 => "000000000000000000000000",
801 => "000000000000000000000000",
802 => "000000000000000000000000",
803 => "000000000000000000000000",
804 => "000000000000000000000000",
805 => "001100110100100110000110",
806 => "010010101000010111101111",
807 => "001011100100101011001100",
808 => "001010100100100011001001",
809 => "010010101000010111101011",
810 => "001110000100110010010100",
811 => "000000000000000000000000",
812 => "000000000000000000000000",
813 => "000000000000000000000000",
814 => "000000000000000000000000",
815 => "000000000000000000000000",
816 => "000000000000000000000000",
817 => "000000000000000000000000",
818 => "000000000000000000000000",
819 => "000000000000000000000000",
820 => "000000000000000000000000",
821 => "000000000000000000000000",
822 => "000000000000000000000000",
823 => "000000000000000000000000",
824 => "000000000000000000000000",
825 => "000000000000000000000000",
826 => "000000010000000000000000",
827 => "000101110001010000010011",
828 => "000000100000001000000010",
829 => "000000000000000000000000",
830 => "000000000000000000000000",
831 => "000000000000000000000000",
832 => "000000000000000000000000",
833 => "000000000000000000000000",
834 => "000000000000000000000000",
835 => "000000000000000000000000",
836 => "000000000000000000000000",
837 => "000000000000000000000000",
838 => "000000000000000000000000",
839 => "000000000000000000000000",
840 => "000000000000000000000000",
841 => "000000000000000000000000",
842 => "000000000000000000000000",
843 => "000000000000000000000000",
844 => "000000000000000000000000",
845 => "000000000000000000000000",
846 => "000000000000000000000000",
847 => "000000000000000000000000",
848 => "000000000000000000000000",
849 => "000000000000000000000000",
850 => "000000000000000000000000",
851 => "000000000000000000000000",
852 => "000000000000000000000000",
853 => "000000000000000000000000",
854 => "000000000000000000000000",
855 => "000000000000000000000000",
856 => "000000000000000000000000",
857 => "000001010000010100000101",
858 => "000110110001100100011001",
859 => "000000000000000000000000",
860 => "000000000000000000000000",
861 => "000000000000000000000000",
862 => "000000000000000000000000",
863 => "000000000000000000000000",
864 => "000000000000000000000000",
865 => "000000000000000000000000",
866 => "000000000000000000000000",
867 => "000000000000000000000000",
868 => "000000000000000000000000",
869 => "000000000000000000000000",
870 => "000000000000000000000000",
871 => "000000000000000000000000",
872 => "000000000000000000000000",
873 => "000000000000000000000000",
874 => "000000000000000000000000",
875 => "001100010100001010001000",
876 => "010010001000001111110001",
877 => "001010000011111111001100",
878 => "001010010011101011001010",
879 => "010010011000001111110001",
880 => "001100100100101010001101",
881 => "000000000000000000000000",
882 => "000000000000000000000000",
883 => "000000000000000000000000",
884 => "000000000000000000000000",
885 => "000000000000000000000000",
886 => "000000000000000000000000",
887 => "000000000000000000000000",
888 => "000000000000000000000000",
889 => "000000000000000000000000",
890 => "000000000000000000000000",
891 => "000000000000000000000000",
892 => "000000000000000000000000",
893 => "000000000000000000000000",
894 => "000000000000000000000000",
895 => "000000000000000000000000",
896 => "000000000000000000000000",
897 => "000110010001100000011000",
898 => "000001100000011000000101",
899 => "000000000000000000000000",
900 => "000000000000000000000000",
901 => "000000000000000000000000",
902 => "000000000000000000000000",
903 => "000000000000000000000000",
904 => "000000000000000000000000",
905 => "000000000000000000000000",
906 => "000000000000000000000000",
907 => "000000000000000000000000",
908 => "000000000000000000000000",
909 => "000000000000000000000000",
910 => "000000000000000000000000",
911 => "000000000000000000000000",
912 => "000000000000000000000000",
913 => "000000000000000000000000",
914 => "000000000000000000000000",
915 => "000000000000000000000000",
916 => "000000000000000000000000",
917 => "000000000000000000000000",
918 => "000000000000000000000000",
919 => "000000000000000000000000",
920 => "000000000000000000000000",
921 => "000000000000000000000000",
922 => "000000000000000000000000",
923 => "000000000000000000000000",
924 => "000000000000000000000000",
925 => "000000000000000000000000",
926 => "000000000000000000000000",
927 => "000011100000111000001100",
928 => "000110000001101000010100",
929 => "000000000000000000000000",
930 => "000000000000000000000000",
931 => "000000000000000000000000",
932 => "000000000000000000000000",
933 => "000000000000000000000000",
934 => "000000000000000000000000",
935 => "000000000000000000000000",
936 => "000000000000000000000000",
937 => "000000000000000000000000",
938 => "000000000000000000000000",
939 => "000000000000000000000000",
940 => "000000000000000000000000",
941 => "000000000000000000000000",
942 => "000000000000000000000000",
943 => "000000000000000000000000",
944 => "000000000000000000000000",
945 => "000011110001010000110000",
946 => "010100110111100111101010",
947 => "001100010011101111010000",
948 => "001010100011110011001011",
949 => "010100110111100111101110",
950 => "000100000001010100101100",
951 => "000000000000000000000000",
952 => "000000000000000000000000",
953 => "000000000000000000000000",
954 => "000000000000000000000000",
955 => "000000000000000000000000",
956 => "000000000000000000000000",
957 => "000000000000000000000000",
958 => "000000000000000000000000",
959 => "000000000000000000000000",
960 => "000000000000000000000000",
961 => "000000000000000000000000",
962 => "000000000000000000000000",
963 => "000000000000000000000000",
964 => "000000000000000000000000",
965 => "000000000000000000000000",
966 => "000000000000000000000000",
967 => "000101110001100000010100",
968 => "000011100000111000001100",
969 => "000000000000000000000000",
970 => "000000000000000000000000",
971 => "000000000000000000000000",
972 => "000000000000000000000000",
973 => "000000000000000000000000",
974 => "000000000000000000000000",
975 => "000000000000000000000000",
976 => "000000000000000000000000",
977 => "000000000000000000000000",
978 => "000000000000000000000000",
979 => "000000000000000000000000",
980 => "000000000000000000000000",
981 => "000000000000000000000000",
982 => "000000000000000000000000",
983 => "000000000000000000000000",
984 => "000000000000000000000000",
985 => "000000000000000000000000",
986 => "000000000000000000000000",
987 => "000000000000000000000000",
988 => "000000000000000000000000",
989 => "000000000000000000000000",
990 => "000000000000000000000000",
991 => "000000000000000000000000",
992 => "000000000000000000000000",
993 => "000000000000000000000000",
994 => "000000000000000000000000",
995 => "000000000000000000000000",
996 => "000000000000000000000000",
997 => "000011100001000000001011",
998 => "000101100001011100010010",
999 => "000000000000000000000000",
1000 => "000000000000000000000000",
1001 => "000000000000000000000000",
1002 => "000000000000000000000000",
1003 => "000000000000000000000000",
1004 => "000000000000000000000000",
1005 => "000000000000000000000000",
1006 => "000000000000000000000000",
1007 => "000000000000000000000000",
1008 => "000000000000000000000000",
1009 => "000000000000000000000000",
1010 => "000000000000000000000000",
1011 => "000000000000000000000000",
1012 => "000000000000000000000000",
1013 => "000000000000000000000000",
1014 => "000000000000000000000000",
1015 => "000000000000000100000010",
1016 => "000100110001111001001100",
1017 => "001001100010101010110000",
1018 => "000111100010100110100111",
1019 => "000100110001111101001101",
1020 => "000000000000000100000010",
1021 => "000000000000000000000000",
1022 => "000000000000000000000000",
1023 => "000000000000000000000000",
1024 => "000000000000000000000000",
1025 => "000000000000000000000000",
1026 => "000000000000000000000000",
1027 => "000000000000000000000000",
1028 => "000000000000000000000000",
1029 => "000000000000000000000000",
1030 => "000000000000000000000000",
1031 => "000000000000000000000000",
1032 => "000000000000000000000000",
1033 => "000000000000000000000000",
1034 => "000000000000000000000000",
1035 => "000000000000000000000000",
1036 => "000000000000000000000000",
1037 => "000101010001010100010010",
1038 => "000011110000111100001100",
1039 => "000000000000000000000000",
1040 => "000000000000000000000000",
1041 => "000000000000000000000000",
1042 => "000000000000000000000000",
1043 => "000000000000000000000000",
1044 => "000000000000000000000000",
1045 => "000000000000000000000000",
1046 => "000000000000000000000000",
1047 => "000000000000000000000000",
1048 => "000000000000000000000000",
1049 => "000000000000000000000000",
1050 => "000000000000000000000000",
1051 => "000000000000000000000000",
1052 => "000000000000000000000000",
1053 => "000000000000000000000000",
1054 => "000000000000000000000000",
1055 => "000000000000000000000000",
1056 => "000000000000000000000000",
1057 => "000000000000000000000000",
1058 => "000000000000000000000000",
1059 => "000000000000000000000000",
1060 => "000000000000000000000000",
1061 => "000000000000000000000000",
1062 => "000000000000000000000000",
1063 => "000000000000000000000000",
1064 => "000000000000000000000000",
1065 => "000000000000000000000000",
1066 => "000000000000000000000000",
1067 => "000110100001101100010111",
1068 => "000010010000100000000110",
1069 => "000000000000000000000000",
1070 => "000000000000000000000000",
1071 => "000000000000000000000000",
1072 => "000000000000000000000000",
1073 => "000000000000000000000000",
1074 => "000000000000000000000000",
1075 => "000000000000000000000000",
1076 => "000000000000000000000000",
1077 => "000000000000000000000000",
1078 => "000000000000000000000000",
1079 => "000000000000000000000000",
1080 => "000000000000000000000000",
1081 => "000000000000000000000000",
1082 => "000000000000000000000000",
1083 => "000000010000000100001100",
1084 => "000100010001001001110011",
1085 => "000100010001001001111001",
1086 => "000000100000001000110011",
1087 => "000000110000001101011101",
1088 => "000001000000010000111110",
1089 => "000000010000000100100010",
1090 => "000011110001000101110000",
1091 => "000100010001001101101101",
1092 => "000000010000000100001011",
1093 => "000000000000000000000000",
1094 => "000000000000000000000000",
1095 => "000000000000000000000000",
1096 => "000000000000000000000000",
1097 => "000000000000000000000000",
1098 => "000000000000000000000000",
1099 => "000000000000000000000000",
1100 => "000000000000000000000000",
1101 => "000000000000000000000000",
1102 => "000000000000000000000000",
1103 => "000000000000000000000000",
1104 => "000000000000000000000000",
1105 => "000000000000000000000000",
1106 => "000000000000000000000000",
1107 => "000010000000100000000110",
1108 => "000110110001101100011001",
1109 => "000000000000000000000000",
1110 => "000000000000000000000000",
1111 => "000000000000000000000000",
1112 => "000000000000000000000000",
1113 => "000000000000000000000000",
1114 => "000000000000000000000000",
1115 => "000000000000000000000000",
1116 => "000000000000000000000000",
1117 => "000000000000000000000000",
1118 => "000000000000000000000000",
1119 => "000000000000000000000000",
1120 => "000000000000000000000000",
1121 => "000000000000000000000000",
1122 => "000000000000000000000000",
1123 => "000000000000000000000000",
1124 => "000000000000000000000000",
1125 => "000000000000000000000000",
1126 => "000000000000000000000000",
1127 => "000000000000000000000000",
1128 => "000000000000000000000000",
1129 => "000000000000000000000000",
1130 => "000000000000000000000000",
1131 => "000000000000000000000000",
1132 => "000000000000000000000000",
1133 => "000000000000000000000000",
1134 => "000000000000000000000000",
1135 => "000000000000000000000000",
1136 => "000000000000000000000000",
1137 => "000110010001101100010111",
1138 => "000010000000011100000110",
1139 => "000000000000000000000000",
1140 => "000000000000000000000000",
1141 => "000000000000000000000000",
1142 => "000000000000000000000000",
1143 => "000000000000000000000000",
1144 => "000000000000000000000000",
1145 => "000000000000000000000000",
1146 => "000000000000000000000000",
1147 => "000000000000000000000000",
1148 => "000000000000000000000000",
1149 => "000000000000000000000000",
1150 => "000000000000000000000000",
1151 => "000000000000000000000000",
1152 => "000000000000000000000000",
1153 => "000010100000110001001011",
1154 => "000100010001011011010001",
1155 => "000100100001010111011000",
1156 => "000100110001011011001001",
1157 => "000001000000010110101100",
1158 => "000001100000011010011100",
1159 => "000100100001011011000001",
1160 => "000100110001010111011001",
1161 => "000100100001011011010000",
1162 => "000011000000101101010011",
1163 => "000000000000000000000000",
1164 => "000000000000000000000000",
1165 => "000000000000000000000000",
1166 => "000000000000000000000000",
1167 => "000000000000000000000000",
1168 => "000000000000000000000000",
1169 => "000000000000000000000000",
1170 => "000000000000000000000000",
1171 => "000000000000000000000000",
1172 => "000000000000000000000000",
1173 => "000000000000000000000000",
1174 => "000000000000000000000000",
1175 => "000000000000000000000000",
1176 => "000000000000000000000000",
1177 => "000001110000011000000110",
1178 => "000110110001110100011001",
1179 => "000000000000000000000000",
1180 => "000000000000000000000000",
1181 => "000000000000000000000000",
1182 => "000000000000000000000000",
1183 => "000000000000000000000000",
1184 => "000000000000000000000000",
1185 => "000000000000000000000000",
1186 => "000000000000000000000000",
1187 => "000000000000000000000000",
1188 => "000000000000000000000000",
1189 => "000000000000000000000000",
1190 => "000000000000000000000000",
1191 => "000000000000000000000000",
1192 => "000000000000000000000000",
1193 => "000000000000000000000000",
1194 => "000000000000000000000000",
1195 => "000000000000000000000000",
1196 => "000000000000000000000000",
1197 => "000000000000000000000000",
1198 => "000000000000000000000000",
1199 => "000000000000000000000000",
1200 => "000000000000000000000000",
1201 => "000000000000000000000000",
1202 => "000000000000000000000000",
1203 => "000000000000000000000000",
1204 => "000000000000000000000000",
1205 => "000000000000000000000000",
1206 => "000000000000000000000000",
1207 => "000101000001011000010010",
1208 => "000001110000011000000110",
1209 => "000000000000000000000000",
1210 => "000000000000000000000000",
1211 => "000000000000000000000000",
1212 => "000000000000000000000000",
1213 => "000000000000000000000000",
1214 => "000000000000000000000000",
1215 => "000000000000000000000000",
1216 => "000000000000000000000000",
1217 => "000000000000000000000000",
1218 => "000000000000000000000000",
1219 => "000000000000000000000000",
1220 => "000000000000000000000000",
1221 => "000000000000000000000000",
1222 => "000000000000000000000000",
1223 => "000001010000001100101100",
1224 => "000101100001001011000001",
1225 => "000101010001010111010010",
1226 => "000101010001010011010110",
1227 => "000001110000010010101101",
1228 => "000010000000001110110101",
1229 => "000101000001010111010001",
1230 => "000100110001010111010011",
1231 => "000101000001011010111110",
1232 => "000001010000010100101011",
1233 => "000000000000000000000000",
1234 => "000000000000000000000000",
1235 => "000000000000000000000000",
1236 => "000000000000000000000000",
1237 => "000000000000000000000000",
1238 => "000000000000000000000000",
1239 => "000000000000000000000000",
1240 => "000000000000000000000000",
1241 => "000000000000000000000000",
1242 => "000000000000000000000000",
1243 => "000000000000000000000000",
1244 => "000000000000000000000000",
1245 => "000000000000000000000000",
1246 => "000000000000000000000000",
1247 => "000001100000011000000101",
1248 => "000101000001011000010010",
1249 => "000000000000000000000000",
1250 => "000000000000000000000000",
1251 => "000000000000000000000000",
1252 => "000000000000000000000000",
1253 => "000000000000000000000000",
1254 => "000000000000000000000000",
1255 => "000000000000000000000000",
1256 => "000000000000000000000000",
1257 => "000000000000000000000000",
1258 => "000000000000000000000000",
1259 => "000000000000000000000000",
1260 => "000000000000000000000000",
1261 => "000000000000000000000000",
1262 => "000000000000000000000000",
1263 => "000000000000000000000000",
1264 => "000000000000000000000000",
1265 => "000000000000000000000000",
1266 => "000000000000000000000000",
1267 => "000000000000000000000000",
1268 => "000000000000000000000000",
1269 => "000000000000000000000000",
1270 => "000000000000000000000000",
1271 => "000000000000000000000000",
1272 => "000000000000000000000000",
1273 => "000000000000000000000000",
1274 => "000000000000000000000000",
1275 => "000000000000000000000000",
1276 => "000000010000000000000001",
1277 => "000101110001100000010101",
1278 => "000001110000011000000110",
1279 => "000000000000000000000000",
1280 => "000000000000000000000000",
1281 => "000000000000000000000000",
1282 => "000000000000000000000000",
1283 => "000000000000000000000000",
1284 => "000000110000001000000010",
1285 => "000000000000000000000000",
1286 => "000000000000000000000000",
1287 => "000000000000000000000000",
1288 => "000000000000000000000000",
1289 => "000000000000000000000000",
1290 => "000000000000000000000000",
1291 => "000000000000000000000000",
1292 => "000000000000000000000000",
1293 => "000000000000000000000001",
1294 => "000000100000001000100010",
1295 => "000011010000111101110100",
1296 => "000100010001010010110111",
1297 => "000000110000100010101011",
1298 => "000000110000011110101011",
1299 => "000100010001010010111011",
1300 => "000011100000111101111011",
1301 => "000000110000000100101100",
1302 => "000000000000000000000000",
1303 => "000000000000000000000000",
1304 => "000000000000000000000000",
1305 => "000000000000000000000000",
1306 => "000000000000000000000000",
1307 => "000000000000000000000000",
1308 => "000000000000000000000000",
1309 => "000000000000000000000000",
1310 => "000000000000000000000000",
1311 => "000000100000001000000010",
1312 => "000000000000000000000000",
1313 => "000000000000000000000000",
1314 => "000000000000000000000000",
1315 => "000000000000000000000000",
1316 => "000000000000000000000000",
1317 => "000001010000011000000101",
1318 => "000101100001100100010100",
1319 => "000000010000000000000000",
1320 => "000000000000000000000000",
1321 => "000000000000000000000000",
1322 => "000000000000000000000000",
1323 => "000000000000000000000000",
1324 => "000000000000000000000000",
1325 => "000000000000000000000000",
1326 => "000000000000000000000000",
1327 => "000000000000000000000000",
1328 => "000000000000000000000000",
1329 => "000000000000000000000000",
1330 => "000000000000000000000000",
1331 => "000000000000000000000000",
1332 => "000000000000000000000000",
1333 => "000000000000000000000000",
1334 => "000000000000000000000000",
1335 => "000000000000000000000000",
1336 => "000000000000000000000000",
1337 => "000000000000000000000000",
1338 => "000000000000000000000000",
1339 => "000000000000000000000000",
1340 => "000000000000000000000000",
1341 => "000000000000000000000000",
1342 => "000000000000000000000000",
1343 => "000000000000000000000000",
1344 => "000000000000000000000000",
1345 => "000000000000000000000000",
1346 => "000000000000000000000000",
1347 => "000110100001101100011000",
1348 => "000010000000011100000110",
1349 => "000000000000000000000000",
1350 => "000000000000000000000000",
1351 => "000000000000000000000000",
1352 => "000000000000000000000000",
1353 => "000001110000011000000110",
1354 => "001001000010000000011001",
1355 => "000001010000010100000100",
1356 => "000000000000000000000000",
1357 => "000000000000000000000000",
1358 => "000000000000000000000000",
1359 => "000000000000000000000000",
1360 => "000000000000000000000000",
1361 => "000000000000000000000000",
1362 => "000000000000000000000000",
1363 => "000000000000000000000000",
1364 => "000000110000001100001110",
1365 => "000010110000101100100001",
1366 => "000001010000010000111011",
1367 => "000001010000001001111001",
1368 => "000001010000001101110110",
1369 => "000000110000010000111101",
1370 => "000010110000101100100001",
1371 => "000001000000001100010000",
1372 => "000000000000000000000000",
1373 => "000000000000000000000000",
1374 => "000000000000000000000000",
1375 => "000000000000000000000000",
1376 => "000000000000000000000000",
1377 => "000000000000000000000000",
1378 => "000000000000000000000000",
1379 => "000000000000000000000000",
1380 => "000001000000001100000011",
1381 => "001000000010000000011010",
1382 => "000001010000010100000100",
1383 => "000000000000000000000000",
1384 => "000000000000000000000000",
1385 => "000000000000000000000000",
1386 => "000000000000000000000000",
1387 => "000001100000011000000110",
1388 => "000110110001110100011000",
1389 => "000000010000000000000000",
1390 => "000000000000000000000000",
1391 => "000000000000000000000000",
1392 => "000000000000000000000000",
1393 => "000000000000000000000000",
1394 => "000000000000000000000000",
1395 => "000000000000000000000000",
1396 => "000000000000000000000000",
1397 => "000000000000000000000000",
1398 => "000000000000000000000000",
1399 => "000000000000000000000000",
1400 => "000000000000000000000000",
1401 => "000000000000000000000000",
1402 => "000000000000000000000000",
1403 => "000000000000000000000000",
1404 => "000000000000000000000000",
1405 => "000000000000000000000000",
1406 => "000000000000000000000000",
1407 => "000000000000000000000000",
1408 => "000000000000000000000000",
1409 => "000000000000000000000000",
1410 => "000000000000000000000000",
1411 => "000000000000000000000000",
1412 => "000000000000000000000000",
1413 => "000000000000000000000000",
1414 => "000000000000000000000000",
1415 => "000000000000000000000000",
1416 => "000000000000000000000000",
1417 => "000110100001101100010111",
1418 => "000001110000011100000111",
1419 => "000000000000000000000000",
1420 => "000000000000000000000000",
1421 => "000000000000000000000000",
1422 => "000000000000000000000000",
1423 => "000101010001010100001110",
1424 => "010100110100101000110100",
1425 => "000011100000110100001000",
1426 => "000000000000000000000000",
1427 => "000000000000000000000000",
1428 => "000000000000000000000000",
1429 => "000000000000000000000000",
1430 => "000000000000000000000000",
1431 => "000000000000000000000000",
1432 => "000000000000000000000000",
1433 => "000010010000100000111011",
1434 => "000111000001110010101010",
1435 => "001010110010111111001101",
1436 => "000010110000110110011111",
1437 => "000000110000011010001010",
1438 => "000000110000010110001101",
1439 => "000011100000110110100101",
1440 => "001011100010111011001101",
1441 => "000110110001110010110101",
1442 => "000010010000100101000101",
1443 => "000000000000000000000000",
1444 => "000000000000000000000000",
1445 => "000000000000000000000000",
1446 => "000000000000000000000000",
1447 => "000000000000000000000000",
1448 => "000000000000000000000000",
1449 => "000000000000000000000000",
1450 => "000011000000100100000111",
1451 => "010100010100101000110100",
1452 => "000100100001000000001101",
1453 => "000000000000000000000000",
1454 => "000000000000000000000000",
1455 => "000000000000000000000000",
1456 => "000000000000000000000000",
1457 => "000001110000011100000110",
1458 => "000110100001110000010111",
1459 => "000000010000000100000001",
1460 => "000000000000000000000000",
1461 => "000000000000000000000000",
1462 => "000000000000000000000000",
1463 => "000000000000000000000000",
1464 => "000000000000000000000000",
1465 => "000000000000000000000000",
1466 => "000000000000000000000000",
1467 => "000000000000000000000000",
1468 => "000000000000000000000000",
1469 => "000000000000000000000000",
1470 => "000000000000000000000000",
1471 => "000000000000000000000000",
1472 => "000000000000000000000000",
1473 => "000000000000000000000000",
1474 => "000000000000000000000000",
1475 => "000000000000000000000000",
1476 => "000000000000000000000000",
1477 => "000000000000000000000000",
1478 => "000000000000000000000000",
1479 => "000000000000000000000000",
1480 => "000000000000000000000000",
1481 => "000000000000000000000000",
1482 => "000000000000000000000000",
1483 => "000000000000000000000000",
1484 => "000000000000000000000000",
1485 => "000000000000000000000000",
1486 => "000000010000000000000000",
1487 => "000101100001011100010011",
1488 => "000001110000011000000110",
1489 => "000000000000000000000000",
1490 => "000000000000000000000000",
1491 => "000000000000000000000000",
1492 => "000000000000000000000000",
1493 => "000100100001000100001001",
1494 => "011001110101110001000011",
1495 => "000100000000111100001001",
1496 => "000000000000000000000000",
1497 => "000000000000000000000000",
1498 => "000000000000000000000000",
1499 => "000000000000000000000000",
1500 => "000000000000000000000000",
1501 => "000000000000000000000000",
1502 => "000000010000000100000101",
1503 => "000101010001011010101111",
1504 => "001100010011011011010000",
1505 => "001101010011101111010010",
1506 => "001000010010001011010100",
1507 => "000010000000100010110111",
1508 => "000010000000100010111010",
1509 => "000111110010001011001111",
1510 => "001101000011101111001111",
1511 => "001101000011100111001101",
1512 => "000101100001011010101111",
1513 => "000000010000000100000101",
1514 => "000000000000000000000000",
1515 => "000000000000000000000000",
1516 => "000000000000000000000000",
1517 => "000000000000000000000000",
1518 => "000000000000000000000000",
1519 => "000000000000000000000000",
1520 => "000011010000101100001000",
1521 => "011001100101100101000000",
1522 => "000011100000110100001001",
1523 => "000000000000000000000000",
1524 => "000000000000000000000000",
1525 => "000000000000000000000000",
1526 => "000000000000000000000000",
1527 => "000001100000011000000101",
1528 => "000101100001100000010100",
1529 => "000000000000000000000000",
1530 => "000000000000000000000000",
1531 => "000000000000000000000000",
1532 => "000000000000000000000000",
1533 => "000000000000000000000000",
1534 => "000000000000000000000000",
1535 => "000000000000000000000000",
1536 => "000000000000000000000000",
1537 => "000000000000000000000000",
1538 => "000000000000000000000000",
1539 => "000000000000000000000000",
1540 => "000000000000000000000000",
1541 => "000000000000000000000000",
1542 => "000000000000000000000000",
1543 => "000000000000000000000000",
1544 => "000000000000000000000000",
1545 => "000000000000000000000000",
1546 => "000000000000000000000000",
1547 => "000000000000000000000000",
1548 => "000000000000000000000000",
1549 => "000000000000000000000000",
1550 => "000000000000000000000000",
1551 => "000000000000000000000000",
1552 => "000000000000000000000000",
1553 => "000000000000000000000000",
1554 => "000000000000000000000000",
1555 => "000000000000000000000000",
1556 => "000000000000000000000000",
1557 => "000101110001100000010100",
1558 => "000001100000011000000101",
1559 => "000000000000000000000000",
1560 => "000000000000000000000000",
1561 => "000000000000000000000000",
1562 => "000000000000000000000000",
1563 => "000000110000001100000010",
1564 => "001001100010000000010111",
1565 => "000011100001000000001101",
1566 => "000000000000000000000000",
1567 => "000000000000000000000000",
1568 => "000000000000000000000000",
1569 => "000000000000000000000000",
1570 => "000000000000000000000000",
1571 => "000000000000000000000000",
1572 => "000000010000000100000101",
1573 => "000101000001011110100010",
1574 => "001011000011001011010000",
1575 => "001110010011111011001111",
1576 => "001000000010001111001000",
1577 => "000010000000100010101111",
1578 => "000001100000100010101001",
1579 => "000111010010000111001101",
1580 => "001110100011111011001110",
1581 => "001011110011001111010000",
1582 => "000110000001011010101010",
1583 => "000000010000000000000100",
1584 => "000000000000000000000000",
1585 => "000000000000000000000000",
1586 => "000000000000000000000000",
1587 => "000000000000000000000000",
1588 => "000000000000000000000000",
1589 => "000000000000000000000000",
1590 => "000011100000110100001011",
1591 => "001001010010001100011000",
1592 => "000000110000001000000010",
1593 => "000000000000000000000000",
1594 => "000000000000000000000000",
1595 => "000000000000000000000000",
1596 => "000000000000000000000000",
1597 => "000001100000011000000101",
1598 => "000101100001100000010100",
1599 => "000000000000000000000000",
1600 => "000000000000000000000000",
1601 => "000000000000000000000000",
1602 => "000000000000000000000000",
1603 => "000000000000000000000000",
1604 => "000000000000000000000000",
1605 => "000000000000000000000000",
1606 => "000000000000000000000000",
1607 => "000000000000000000000000",
1608 => "000000000000000000000000",
1609 => "000000000000000000000000",
1610 => "000000000000000000000000",
1611 => "000000000000000000000000",
1612 => "000000000000000000000000",
1613 => "000000000000000000000000",
1614 => "000000000000000000000000",
1615 => "000000000000000000000000",
1616 => "000000000000000000000000",
1617 => "000000000000000000000000",
1618 => "000000000000000000000000",
1619 => "000000000000000000000000",
1620 => "000000000000000000000000",
1621 => "000000000000000000000000",
1622 => "000000000000000000000000",
1623 => "000000000000000000000000",
1624 => "000000000000000000000000",
1625 => "000000000000000000000000",
1626 => "000000010000000100000001",
1627 => "000110100001110100011010",
1628 => "000001110000011000000110",
1629 => "000000000000000000000000",
1630 => "000000000000000000000000",
1631 => "000000000000000000000000",
1632 => "000000000000000000000000",
1633 => "000000000000000000000000",
1634 => "000001010000001100000100",
1635 => "000111000001100100011001",
1636 => "000001010000010000000011",
1637 => "000000000000000000000000",
1638 => "000000000000000000000000",
1639 => "000000000000000000000000",
1640 => "000000000000000000000000",
1641 => "000000000000000000000000",
1642 => "000000000000000000000000",
1643 => "000001010000010000100101",
1644 => "000101010001010010010111",
1645 => "001001100010110110101111",
1646 => "000010100000110110000001",
1647 => "000000100000001100111111",
1648 => "000000110000001100111011",
1649 => "000010110000110110000101",
1650 => "001010100010110110101111",
1651 => "000100100001100010011100",
1652 => "000001100000010000110001",
1653 => "000000000000000000000000",
1654 => "000000000000000000000000",
1655 => "000000000000000000000000",
1656 => "000000000000000000000000",
1657 => "000000000000000000000000",
1658 => "000000000000000000000000",
1659 => "000000110000001100000010",
1660 => "000110010001100100010101",
1661 => "000001010000010000000100",
1662 => "000000000000000000000000",
1663 => "000000000000000000000000",
1664 => "000000000000000000000000",
1665 => "000000000000000000000000",
1666 => "000000000000000000000000",
1667 => "000001100000011100000101",
1668 => "000110000001110100011000",
1669 => "000000010000000000000000",
1670 => "000000000000000000000000",
1671 => "000000000000000000000000",
1672 => "000000000000000000000000",
1673 => "000000000000000000000000",
1674 => "000000000000000000000000",
1675 => "000000000000000000000000",
1676 => "000000000000000000000000",
1677 => "000000000000000000000000",
1678 => "000000000000000000000000",
1679 => "000000000000000000000000",
1680 => "000000000000000000000000",
1681 => "000000000000000000000000",
1682 => "000000000000000000000000",
1683 => "000000000000000000000000",
1684 => "000000000000000000000000",
1685 => "000000000000000000000000",
1686 => "000000000000000000000000",
1687 => "000000000000000000000000",
1688 => "000000000000000000000000",
1689 => "000000000000000000000000",
1690 => "000000000000000000000000",
1691 => "000000000000000000000000",
1692 => "000000000000000000000000",
1693 => "000000000000000000000000",
1694 => "000000000000000000000000",
1695 => "000000000000000000000000",
1696 => "000000010000000100000001",
1697 => "000111000001111000011011",
1698 => "000010000000011000000111",
1699 => "000000000000000000000000",
1700 => "000000000000000000000000",
1701 => "000000000000000000000000",
1702 => "000000000000000000000000",
1703 => "000000000000000000000000",
1704 => "000000000000000000000000",
1705 => "000110000001010000010001",
1706 => "000110000001010100010001",
1707 => "000000000000000000000000",
1708 => "000000000000000000000000",
1709 => "000000000000000000000000",
1710 => "000000000000000000000000",
1711 => "000000000000000000000000",
1712 => "000000000000000000000000",
1713 => "000000000000000000000000",
1714 => "000000100000000100000111",
1715 => "000001110000011100100110",
1716 => "000001110000011100111100",
1717 => "000000110000010000011101",
1718 => "000001000000001100011100",
1719 => "000001110000100000111101",
1720 => "000001110000100000100111",
1721 => "000000010000001000001001",
1722 => "000000000000000000000000",
1723 => "000000000000000000000000",
1724 => "000000000000000000000000",
1725 => "000000000000000000000000",
1726 => "000000000000000000000000",
1727 => "000000000000000000000000",
1728 => "000000000000000000000000",
1729 => "000101100001001100010000",
1730 => "000110000001011000010011",
1731 => "000000000000000000000000",
1732 => "000000000000000000000000",
1733 => "000000000000000000000000",
1734 => "000000000000000000000000",
1735 => "000000000000000000000000",
1736 => "000000000000000000000000",
1737 => "000001110000011000000110",
1738 => "000111000001111000011010",
1739 => "000000010000000000000000",
1740 => "000000000000000000000000",
1741 => "000000000000000000000000",
1742 => "000000000000000000000000",
1743 => "000000000000000000000000",
1744 => "000000000000000000000000",
1745 => "000000000000000000000000",
1746 => "000000000000000000000000",
1747 => "000000000000000000000000",
1748 => "000000000000000000000000",
1749 => "000000000000000000000000",
1750 => "000000000000000000000000",
1751 => "000000000000000000000000",
1752 => "000000000000000000000000",
1753 => "000000000000000000000000",
1754 => "000000000000000000000000",
1755 => "000000000000000000000000",
1756 => "000000000000000000000000",
1757 => "000000000000000000000000",
1758 => "000000000000000000000000",
1759 => "000000000000000000000000",
1760 => "000000000000000000000000",
1761 => "000000000000000000000000",
1762 => "000000000000000000000000",
1763 => "000000000000000000000000",
1764 => "000000000000000000000000",
1765 => "000000000000000000000000",
1766 => "000000010000000000000001",
1767 => "000110000001101000010111",
1768 => "000001110000011000000101",
1769 => "000000000000000000000000",
1770 => "000000000000000000000000",
1771 => "000000000000000000000000",
1772 => "000000000000000000000000",
1773 => "000000000000000000000000",
1774 => "000000000000000000000000",
1775 => "000100100000111100001101",
1776 => "001001110010010000011100",
1777 => "000000000000000000000000",
1778 => "000000000000000000000000",
1779 => "000000000000000000000000",
1780 => "000000000000000000000000",
1781 => "000000000000000000000000",
1782 => "000000000000000000000000",
1783 => "000000110000001100001011",
1784 => "010001110101100010011001",
1785 => "010011010111001011011101",
1786 => "010010010110001011100000",
1787 => "000011010001000010000011",
1788 => "000011010000111101111100",
1789 => "010010100110000111011110",
1790 => "010011000111001011011101",
1791 => "010010110110001110100110",
1792 => "000000110000010100010010",
1793 => "000000000000000000000000",
1794 => "000000000000000000000000",
1795 => "000000000000000000000000",
1796 => "000000000000000000000000",
1797 => "000000000000000000000000",
1798 => "000000000000000000000000",
1799 => "001000100010000000011100",
1800 => "000100100001000100001111",
1801 => "000000000000000000000000",
1802 => "000000000000000000000000",
1803 => "000000000000000000000000",
1804 => "000000000000000000000000",
1805 => "000000000000000000000000",
1806 => "000000000000000000000000",
1807 => "000001100000011000000101",
1808 => "000110000001101000010110",
1809 => "000000010000000000000001",
1810 => "000000000000000000000000",
1811 => "000000000000000000000000",
1812 => "000000000000000000000000",
1813 => "000000000000000000000000",
1814 => "000000000000000000000000",
1815 => "000000000000000000000000",
1816 => "000000000000000000000000",
1817 => "000000000000000000000000",
1818 => "000000000000000000000000",
1819 => "000000000000000000000000",
1820 => "000000000000000000000000",
1821 => "000000000000000000000000",
1822 => "000000000000000000000000",
1823 => "000000000000000000000000",
1824 => "000000000000000000000000",
1825 => "000000000000000000000000",
1826 => "000000000000000000000000",
1827 => "000000000000000000000000",
1828 => "000000000000000000000000",
1829 => "000000000000000000000000",
1830 => "000000000000000000000000",
1831 => "000000000000000000000000",
1832 => "000000000000000000000000",
1833 => "000000000000000000000000",
1834 => "000000000000000000000000",
1835 => "000000000000000000000000",
1836 => "000000010000000100000001",
1837 => "000111100010001000011101",
1838 => "000001100000011000000101",
1839 => "000000000000000000000000",
1840 => "000000000000000000000000",
1841 => "000000000000000000000000",
1842 => "000000000000000000000000",
1843 => "000000000000000000000000",
1844 => "000000000000000000000000",
1845 => "000011000000101100001000",
1846 => "001010110010100100011011",
1847 => "000001010000001100000011",
1848 => "000000000000000000000000",
1849 => "000000000000000000000000",
1850 => "000000000000000000000000",
1851 => "000000000000000000000000",
1852 => "000000000000000000000001",
1853 => "001001000010110101100110",
1854 => "010110011000110111101110",
1855 => "010001101000110011110100",
1856 => "010001100111001111110001",
1857 => "000011010001000110100100",
1858 => "000010110001000010011110",
1859 => "010001100111001111101110",
1860 => "010010011000101011110101",
1861 => "010110011000111011110010",
1862 => "001011100011100010000110",
1863 => "000000000000000000000000",
1864 => "000000000000000000000000",
1865 => "000000000000000000000000",
1866 => "000000000000000000000000",
1867 => "000000000000000000000000",
1868 => "000000110000001000000010",
1869 => "001001110010010100011101",
1870 => "000011000000101100001001",
1871 => "000000000000000000000000",
1872 => "000000000000000000000000",
1873 => "000000000000000000000000",
1874 => "000000000000000000000000",
1875 => "000000000000000000000000",
1876 => "000000000000000000000000",
1877 => "000001010000011000000101",
1878 => "000111100010001000011101",
1879 => "000000010000000100000001",
1880 => "000000000000000000000000",
1881 => "000000000000000000000000",
1882 => "000000000000000000000000",
1883 => "000000000000000000000000",
1884 => "000000000000000000000000",
1885 => "000000000000000000000000",
1886 => "000000000000000000000000",
1887 => "000000000000000000000000",
1888 => "000000000000000000000000",
1889 => "000000000000000000000000",
1890 => "000000000000000000000000",
1891 => "000000000000000000000000",
1892 => "000000000000000000000000",
1893 => "000000000000000000000000",
1894 => "000000000000000000000000",
1895 => "000000000000000000000000",
1896 => "000000000000000000000000",
1897 => "000000000000000000000000",
1898 => "000000000000000000000000",
1899 => "000000000000000000000000",
1900 => "000000000000000000000000",
1901 => "000000000000000000000000",
1902 => "000000000000000000000000",
1903 => "000000000000000000000000",
1904 => "000000000000000000000000",
1905 => "000000000000000000000000",
1906 => "000000010000000100000001",
1907 => "001010000011001000101011",
1908 => "000001100000011100000110",
1909 => "000000000000000000000000",
1910 => "000000000000000000000000",
1911 => "000000000000000000000000",
1912 => "000000000000000000000000",
1913 => "000000000000000000000000",
1914 => "000000000000000000000000",
1915 => "000100100000111100001100",
1916 => "011011010110010001001001",
1917 => "000011100000110000001001",
1918 => "000000000000000000000000",
1919 => "000000000000000000000100",
1920 => "000000110000000100010010",
1921 => "000000000000000000000000",
1922 => "000000110000001100000110",
1923 => "010100010110110011001110",
1924 => "010011111000111011110100",
1925 => "010010101000000011101111",
1926 => "001111110101000111000100",
1927 => "000011110000110101001000",
1928 => "000010100000110001000111",
1929 => "010000010100111111000100",
1930 => "010010001000000111101101",
1931 => "010010001001000011110000",
1932 => "010100010111001011010011",
1933 => "000000110000001100000110",
1934 => "000000000000000000000001",
1935 => "000001000000000100010111",
1936 => "000000010000000000000101",
1937 => "000000000000000000000000",
1938 => "000011000000101100001000",
1939 => "011010100110001001000101",
1940 => "000100100001000000001101",
1941 => "000000000000000000000000",
1942 => "000000000000000000000000",
1943 => "000000000000000000000000",
1944 => "000000000000000000000000",
1945 => "000000000000000000000000",
1946 => "000000000000000000000000",
1947 => "000001110000011100000110",
1948 => "001011000011000000101100",
1949 => "000000010000000100000001",
1950 => "000000000000000000000000",
1951 => "000000000000000000000000",
1952 => "000000000000000000000000",
1953 => "000000000000000000000000",
1954 => "000000000000000000000000",
1955 => "000000000000000000000000",
1956 => "000000000000000000000000",
1957 => "000000000000000000000000",
1958 => "000000000000000000000000",
1959 => "000000000000000000000000",
1960 => "000000000000000000000000",
1961 => "000000000000000000000000",
1962 => "000000000000000000000000",
1963 => "000000000000000000000000",
1964 => "000000000000000000000000",
1965 => "000000000000000000000000",
1966 => "000000000000000000000000",
1967 => "000000000000000000000000",
1968 => "000000000000000000000000",
1969 => "000000000000000000000000",
1970 => "000000000000000000000000",
1971 => "000000000000000000000000",
1972 => "000000000000000000000000",
1973 => "000000000000000000000000",
1974 => "000000000000000000000000",
1975 => "000000000000000000000000",
1976 => "000000010000000100000001",
1977 => "000100110001101000010100",
1978 => "000001010000010100000101",
1979 => "000000000000000000000000",
1980 => "000000000000000000000000",
1981 => "000000000000000000000000",
1982 => "000000000000000000000000",
1983 => "000000000000000000000000",
1984 => "000000000000000000000000",
1985 => "000000000000000000000000",
1986 => "001100110010110100011111",
1987 => "000011100000111000001001",
1988 => "000000010000000100001000",
1989 => "000001110000010101011100",
1990 => "000001100000010101100000",
1991 => "000001000000001100101001",
1992 => "000000110000001100000110",
1993 => "010010100101011010101010",
1994 => "010000000101010110110101",
1995 => "001101110100011010000010",
1996 => "000011010000111000110011",
1997 => "000000010000010000010000",
1998 => "000000110000001100001101",
1999 => "000011010000110000110100",
2000 => "001101110100011010000000",
2001 => "010000110100111110111000",
2002 => "010010010101100110110011",
2003 => "000000100000001100000101",
2004 => "000001010000000100100101",
2005 => "000010010000010101100000",
2006 => "000010010000011001010100",
2007 => "000000010000000000000110",
2008 => "000011100000110100001000",
2009 => "001101000010111000011100",
2010 => "000000000000000000000000",
2011 => "000000000000000000000000",
2012 => "000000000000000000000000",
2013 => "000000000000000000000000",
2014 => "000000000000000000000000",
2015 => "000000000000000000000000",
2016 => "000000000000000000000000",
2017 => "000001000000010100000100",
2018 => "000101000001100100010100",
2019 => "000000010000000100000001",
2020 => "000000000000000000000000",
2021 => "000000000000000000000000",
2022 => "000000000000000000000000",
2023 => "000000000000000000000000",
2024 => "000000000000000000000000",
2025 => "000000000000000000000000",
2026 => "000000000000000000000000",
2027 => "000000000000000000000000",
2028 => "000000000000000000000000",
2029 => "000000000000000000000000",
2030 => "000000000000000000000000",
2031 => "000000000000000000000000",
2032 => "000000000000000000000000",
2033 => "000000000000000000000000",
2034 => "000000000000000000000000",
2035 => "000000000000000000000000",
2036 => "000000000000000000000000",
2037 => "000000000000000000000000",
2038 => "000000000000000000000000",
2039 => "000000000000000000000000",
2040 => "000000000000000000000000",
2041 => "000000000000000000000000",
2042 => "000000000000000000000000",
2043 => "000000000000000000000000",
2044 => "000000000000000000000000",
2045 => "000000000000000000000000",
2046 => "000000010000000100000001",
2047 => "001010110011010000101101",
2048 => "000001100000011000000101",
2049 => "000000000000000000000000",
2050 => "000000000000000000000000",
2051 => "000000000000000000000000",
2052 => "000000000000000000000000",
2053 => "000000000000000000000000",
2054 => "000000110000001000000010",
2055 => "000000100000000100000001",
2056 => "010111010101010100111100",
2057 => "001110000011010100100010",
2058 => "000000010000000100000111",
2059 => "000001000000010100111110",
2060 => "000001110000001101011000",
2061 => "000001010000010101001000",
2062 => "000000000000000000000010",
2063 => "000000000000000000000100",
2064 => "000001100000011001000100",
2065 => "000001110000011101111000",
2066 => "000001100000100101111011",
2067 => "000001000000001101000011",
2068 => "000001100000001001001000",
2069 => "000010000000011101111001",
2070 => "000010010000011101110101",
2071 => "000010010000011001010110",
2072 => "000000100000001000001101",
2073 => "000000000000000000000001",
2074 => "000001110000010001000010",
2075 => "000001100000010001011001",
2076 => "000001010000001101000000",
2077 => "000000100000000100001011",
2078 => "001101000011000000100000",
2079 => "010111100101011000111110",
2080 => "000000010000000100000001",
2081 => "000000100000001000000010",
2082 => "000000000000000000000000",
2083 => "000000000000000000000000",
2084 => "000000000000000000000000",
2085 => "000000000000000000000000",
2086 => "000000000000000000000000",
2087 => "000001100000011000000101",
2088 => "001011110011001000101110",
2089 => "000000100000001000000010",
2090 => "000000000000000000000000",
2091 => "000000000000000000000000",
2092 => "000000000000000000000000",
2093 => "000000000000000000000000",
2094 => "000000000000000000000000",
2095 => "000000000000000000000000",
2096 => "000000000000000000000000",
2097 => "000000000000000000000000",
2098 => "000000000000000000000000",
2099 => "000000000000000000000000",
2100 => "000000000000000000000000",
2101 => "000000000000000000000000",
2102 => "000000000000000000000000",
2103 => "000000000000000000000000",
2104 => "000000000000000000000000",
2105 => "000000000000000000000000",
2106 => "000000000000000000000000",
2107 => "000000000000000000000000",
2108 => "000000000000000000000000",
2109 => "000000000000000000000000",
2110 => "000000000000000000000000",
2111 => "000000000000000000000000",
2112 => "000000000000000000000000",
2113 => "000000000000000000000000",
2114 => "000000000000000000000000",
2115 => "000000000000000000000000",
2116 => "000000010000000000000001",
2117 => "000111110010010100100000",
2118 => "000110000001101100011001",
2119 => "000000000000000000000000",
2120 => "000000000000000000000000",
2121 => "000000000000000000000000",
2122 => "000000000000000000000000",
2123 => "000000100000000100000010",
2124 => "000110000001010000010101",
2125 => "000011110000111000001001",
2126 => "010000110100000000100100",
2127 => "010010000100001000101101",
2128 => "000001000000010000001000",
2129 => "000000110000001000101001",
2130 => "000001000000001000111111",
2131 => "000001100000010101001000",
2132 => "000000000000000000000010",
2133 => "000001100000011100111100",
2134 => "000011110001001011000100",
2135 => "000011110001001011001010",
2136 => "000011100001001011001100",
2137 => "000001110000010010011010",
2138 => "000001000000010110010101",
2139 => "000100000001000111001000",
2140 => "000011110001000111001100",
2141 => "000100000001001111000100",
2142 => "000010100000011101001010",
2143 => "000000000000000000000001",
2144 => "000010000000010001000000",
2145 => "000000110000001101000010",
2146 => "000000110000001100100110",
2147 => "000001100000010100001101",
2148 => "010001100011111100101011",
2149 => "010000100100001000100110",
2150 => "000011010000110000001001",
2151 => "000101010001010100010010",
2152 => "000000010000000100000001",
2153 => "000000000000000000000000",
2154 => "000000000000000000000000",
2155 => "000000000000000000000000",
2156 => "000000000000000000000000",
2157 => "000101010001101000010110",
2158 => "000111010010010100100000",
2159 => "000000000000000000000000",
2160 => "000000000000000000000000",
2161 => "000000000000000000000000",
2162 => "000000000000000000000000",
2163 => "000000000000000000000000",
2164 => "000000000000000000000000",
2165 => "000000000000000000000000",
2166 => "000000000000000000000000",
2167 => "000000000000000000000000",
2168 => "000000000000000000000000",
2169 => "000000000000000000000000",
2170 => "000000000000000000000000",
2171 => "000000000000000000000000",
2172 => "000000000000000000000000",
2173 => "000000000000000000000000",
2174 => "000000000000000000000000",
2175 => "000000000000000000000000",
2176 => "000000000000000000000000",
2177 => "000000000000000000000000",
2178 => "000000000000000000000000",
2179 => "000000000000000000000000",
2180 => "000000000000000000000000",
2181 => "000000000000000000000000",
2182 => "000000000000000000000000",
2183 => "000000000000000000000000",
2184 => "000000000000000000000000",
2185 => "000000000000000000000000",
2186 => "000000010000000000000001",
2187 => "000101100001101100010111",
2188 => "000101110001101100011001",
2189 => "000000000000000000000000",
2190 => "000000000000000000000000",
2191 => "000000000000000000000000",
2192 => "000000000000000000000000",
2193 => "000001000000001100000011",
2194 => "000111110010001100100011",
2195 => "001000110010100000110011",
2196 => "010101010101010100110111",
2197 => "010101110100111000110110",
2198 => "000101010001100000011010",
2199 => "000001100000010001010000",
2200 => "000001010000001101000111",
2201 => "000000110000010000111000",
2202 => "000001000000001100101001",
2203 => "000011100000111110100100",
2204 => "000011110001000111001110",
2205 => "000011110001000111001101",
2206 => "000100000001000111001001",
2207 => "000001010000011001110011",
2208 => "000001000000011101101011",
2209 => "000100010001000111001011",
2210 => "000011110001000011001101",
2211 => "000011100001000111010010",
2212 => "000100000001000010101011",
2213 => "000001000000001000101000",
2214 => "000001010000001000111001",
2215 => "000001000000010001001001",
2216 => "000001010000010001001111",
2217 => "000100110001001100011110",
2218 => "010101110100101100101111",
2219 => "010110110101010000111001",
2220 => "001000010010101100110010",
2221 => "000111010010001100100011",
2222 => "000000110000001100000011",
2223 => "000000000000000000000000",
2224 => "000000000000000000000000",
2225 => "000000000000000000000000",
2226 => "000000000000000000000000",
2227 => "000101110001101100010111",
2228 => "000110000001101100010111",
2229 => "000000000000000000000000",
2230 => "000000000000000000000000",
2231 => "000000000000000000000000",
2232 => "000000000000000000000000",
2233 => "000000000000000000000000",
2234 => "000000000000000000000000",
2235 => "000000000000000000000000",
2236 => "000000000000000000000000",
2237 => "000000000000000000000000",
2238 => "000000000000000000000000",
2239 => "000000000000000000000000",
2240 => "000000000000000000000000",
2241 => "000000000000000000000000",
2242 => "000000000000000000000000",
2243 => "000000000000000000000000",
2244 => "000000000000000000000000",
2245 => "000000000000000000000000",
2246 => "000000000000000000000000",
2247 => "000000000000000000000000",
2248 => "000000000000000000000000",
2249 => "000000000000000000000000",
2250 => "000000000000000000000000",
2251 => "000000000000000000000000",
2252 => "000000000000000000000000",
2253 => "000000000000000000000000",
2254 => "000000000000000000000000",
2255 => "000000000000000000000000",
2256 => "000000010000000100000001",
2257 => "001100000011100100110011",
2258 => "000101110001111100011011",
2259 => "000000000000000000000000",
2260 => "000000000000000000000000",
2261 => "000000000000000000000000",
2262 => "000000000000000000000000",
2263 => "000000100000001000000010",
2264 => "000101110001100100101101",
2265 => "001001010010011101001110",
2266 => "010111100101110000111101",
2267 => "011111100110110100111111",
2268 => "001000010001101100011100",
2269 => "000001000000001100111110",
2270 => "000001010000001101010001",
2271 => "000001000000001101000111",
2272 => "000001100000010001001101",
2273 => "000100100001000110110001",
2274 => "000011110001001111001010",
2275 => "000100010001001010111001",
2276 => "000010000000100101110011",
2277 => "000001000000001100011111",
2278 => "000000100000001000100010",
2279 => "000010000000100101110000",
2280 => "000100010001001010111010",
2281 => "000100010001000111000110",
2282 => "000100010001000110110110",
2283 => "000001100000010001001100",
2284 => "000001100000001001001010",
2285 => "000001010000001101010001",
2286 => "000001010000001101000101",
2287 => "000110000001100100010000",
2288 => "011101000110111001000010",
2289 => "011000100110000100111100",
2290 => "001001000010101001010010",
2291 => "000101110001101000101010",
2292 => "000000100000000100000001",
2293 => "000000000000000000000000",
2294 => "000000000000000000000000",
2295 => "000000000000000000000000",
2296 => "000000000000000000000000",
2297 => "000101100001111000011000",
2298 => "001011110011101000110011",
2299 => "000000010000000100000001",
2300 => "000000000000000000000000",
2301 => "000000000000000000000000",
2302 => "000000000000000000000000",
2303 => "000000000000000000000000",
2304 => "000000000000000000000000",
2305 => "000000000000000000000000",
2306 => "000000000000000000000000",
2307 => "000000000000000000000000",
2308 => "000000000000000000000000",
2309 => "000000000000000000000000",
2310 => "000000000000000000000000",
2311 => "000000000000000000000000",
2312 => "000000000000000000000000",
2313 => "000000000000000000000000",
2314 => "000000000000000000000000",
2315 => "000000000000000000000000",
2316 => "000000000000000000000000",
2317 => "000000000000000000000000",
2318 => "000000000000000000000000",
2319 => "000000000000000000000000",
2320 => "000000000000000000000000",
2321 => "000000000000000000000000",
2322 => "000000000000000000000000",
2323 => "000000000000000000000000",
2324 => "000000000000000000000000",
2325 => "000000000000000000000000",
2326 => "000000000000000000000000",
2327 => "000101010001101100010111",
2328 => "000101110001101100011000",
2329 => "000000000000000000000000",
2330 => "000000000000000000000000",
2331 => "000000000000000000000000",
2332 => "000000000000000000000000",
2333 => "000000100000001000000001",
2334 => "001010010010011100011011",
2335 => "010011000100100001010011",
2336 => "001000100010010101001110",
2337 => "001000110010100000101101",
2338 => "000011010000101000010011",
2339 => "000001100000010001000110",
2340 => "000000110000001101001111",
2341 => "000001010000001101010001",
2342 => "000000110000001000100101",
2343 => "000001110000001101000111",
2344 => "000001100000001101010001",
2345 => "000001000000001100111010",
2346 => "000001000000011000110010",
2347 => "000001000000001000100011",
2348 => "000000110000001100100100",
2349 => "000001100000010100110000",
2350 => "000001000000010000111011",
2351 => "000001000000010101001100",
2352 => "000001100000010001001001",
2353 => "000000100000001000100010",
2354 => "000001000000001101010000",
2355 => "000000110000001101010011",
2356 => "000001100000010101001000",
2357 => "000010110000100100010011",
2358 => "001001000010011000101001",
2359 => "001000110010011001010001",
2360 => "010011000100010001010000",
2361 => "001010100010100000100010",
2362 => "000000110000001000000010",
2363 => "000000000000000000000000",
2364 => "000000000000000000000000",
2365 => "000000000000000000000000",
2366 => "000000000000000000000000",
2367 => "000101110001101100010111",
2368 => "000101110001110000011000",
2369 => "000000000000000000000000",
2370 => "000000000000000000000000",
2371 => "000000000000000000000000",
2372 => "000000000000000000000000",
2373 => "000000000000000000000000",
2374 => "000000000000000000000000",
2375 => "000000000000000000000000",
2376 => "000000000000000000000000",
2377 => "000000000000000000000000",
2378 => "000000000000000000000000",
2379 => "000000000000000000000000",
2380 => "000000000000000000000000",
2381 => "000000000000000000000000",
2382 => "000000000000000000000000",
2383 => "000000000000000000000000",
2384 => "000000000000000000000000",
2385 => "000000000000000000000000",
2386 => "000000000000000000000000",
2387 => "000000000000000000000000",
2388 => "000000000000000000000000",
2389 => "000000000000000000000000",
2390 => "000000000000000000000000",
2391 => "000000000000000000000000",
2392 => "000000000000000000000000",
2393 => "000000000000000000000000",
2394 => "000000000000000000000000",
2395 => "000000000000000000000000",
2396 => "000000010000000100000001",
2397 => "001001100011000000101010",
2398 => "001000010010100000100101",
2399 => "000000000000000000000000",
2400 => "000000000000000000000000",
2401 => "000000000000000000000000",
2402 => "000000000000000000000000",
2403 => "000001010000010000000100",
2404 => "001101100011000100100001",
2405 => "100001010111011101000110",
2406 => "010001100100011101000100",
2407 => "001110010011100000111100",
2408 => "000100100001010100110111",
2409 => "000001000000001000101111",
2410 => "000001000000001001001001",
2411 => "000001000000001101010011",
2412 => "000001000000001100011101",
2413 => "000010010000101100100110",
2414 => "010001110110000010101000",
2415 => "010010000110011011010110",
2416 => "010000110101100111011101",
2417 => "000011100000110110101000",
2418 => "000010100000111010100101",
2419 => "010001000101011111011101",
2420 => "010001110110010111010100",
2421 => "010011000110000110101010",
2422 => "000010110000101100101111",
2423 => "000000100000001100100000",
2424 => "000001010000001101010001",
2425 => "000001010000001101000110",
2426 => "000000100000001100101110",
2427 => "000100010001000100111100",
2428 => "001101000011011000111010",
2429 => "010001110100101001000101",
2430 => "100000100111011001000100",
2431 => "001101100011000100100000",
2432 => "000001000000001100000011",
2433 => "000000000000000000000000",
2434 => "000000000000000000000000",
2435 => "000000000000000000000000",
2436 => "000000000000000000000000",
2437 => "000111110010011100100001",
2438 => "001001110011000100101010",
2439 => "000000010000000100000001",
2440 => "000000000000000000000000",
2441 => "000000000000000000000000",
2442 => "000000000000000000000000",
2443 => "000000000000000000000000",
2444 => "000000000000000000000000",
2445 => "000000000000000000000000",
2446 => "000000000000000000000000",
2447 => "000000000000000000000000",
2448 => "000000000000000000000000",
2449 => "000000000000000000000000",
2450 => "000000000000000000000000",
2451 => "000000000000000000000000",
2452 => "000000000000000000000000",
2453 => "000000000000000000000000",
2454 => "000000000000000000000000",
2455 => "000000000000000000000000",
2456 => "000000000000000000000000",
2457 => "000000000000000000000000",
2458 => "000000000000000000000000",
2459 => "000000000000000000000000",
2460 => "000000000000000000000000",
2461 => "000000000000000000000000",
2462 => "000000000000000000000000",
2463 => "000000000000000000000000",
2464 => "000000000000000000000000",
2465 => "000000000000000000000000",
2466 => "000000000000000000000000",
2467 => "000100010001011100010011",
2468 => "000111000010001100011111",
2469 => "000000000000000000000000",
2470 => "000000000000000000000000",
2471 => "000000000000000000000000",
2472 => "000000000000000000000000",
2473 => "000001110000001100000111",
2474 => "001011000010010100010010",
2475 => "100001110111100101000110",
2476 => "010111110110001000111011",
2477 => "100000100111000101000010",
2478 => "000111110001111000111110",
2479 => "000001100000001100111111",
2480 => "000001010000010101011100",
2481 => "000001000000010101001000",
2482 => "000001000000001000100110",
2483 => "001010010011001010001010",
2484 => "010101011000011011110000",
2485 => "010000111000100111110001",
2486 => "010000100111000011101111",
2487 => "000011000001000010110010",
2488 => "000011000000110110110011",
2489 => "010000100111001111101110",
2490 => "010001001000100111110011",
2491 => "010100111000101011110001",
2492 => "001011110011101010010000",
2493 => "000001010000001000100111",
2494 => "000000110000010001001000",
2495 => "000001110000010001011111",
2496 => "000001100000010000111101",
2497 => "000111110001101100111000",
2498 => "011111100110111001000010",
2499 => "011001110110001000111111",
2500 => "100001110111011001000011",
2501 => "001011010010011100011010",
2502 => "000001000000001000000011",
2503 => "000000000000000000000000",
2504 => "000000000000000000000000",
2505 => "000000000000000000000000",
2506 => "000000000000000000000000",
2507 => "000111010001111100011011",
2508 => "000101010001010100010010",
2509 => "000000000000000000000000",
2510 => "000000000000000000000000",
2511 => "000000000000000000000000",
2512 => "000000000000000000000000",
2513 => "000000000000000000000000",
2514 => "000000000000000000000000",
2515 => "000000000000000000000000",
2516 => "000000000000000000000000",
2517 => "000000000000000000000000",
2518 => "000000000000000000000000",
2519 => "000000000000000000000000",
2520 => "000000000000000000000000",
2521 => "000000000000000000000000",
2522 => "000000000000000000000000",
2523 => "000000000000000000000000",
2524 => "000000000000000000000000",
2525 => "000000000000000000000000",
2526 => "000000000000000000000000",
2527 => "000000000000000000000000",
2528 => "000000000000000000000000",
2529 => "000000000000000000000000",
2530 => "000000000000000000000000",
2531 => "000000000000000000000000",
2532 => "000000000000000000000000",
2533 => "000000000000000000000000",
2534 => "000000000000000000000000",
2535 => "000000000000000000000000",
2536 => "000000000000000000000000",
2537 => "000110100001111000011011",
2538 => "001011000011001100110000",
2539 => "000000110000001100000011",
2540 => "000000000000000000000000",
2541 => "000000000000000000000000",
2542 => "000000000000000000000000",
2543 => "000101010000110000001010",
2544 => "010000110010111100011010",
2545 => "100010010111101001000101",
2546 => "011001000110011001000000",
2547 => "011011110110101100111011",
2548 => "001111010010011000100000",
2549 => "000100000000101000100000",
2550 => "000000110000001000100011",
2551 => "000001010000001101010010",
2552 => "000001110000100101100110",
2553 => "010011110110101011010000",
2554 => "010011101000110011101110",
2555 => "010010100111111111110001",
2556 => "001101110100110111000011",
2557 => "000010110000101101101101",
2558 => "000011000000101001110111",
2559 => "001101110100111011000110",
2560 => "010010001000000111110000",
2561 => "010010011000111011110001",
2562 => "010011110110111111010011",
2563 => "000010100000100101100110",
2564 => "000000110000010001010011",
2565 => "000000110000001000100100",
2566 => "000011100000100000100000",
2567 => "001110100010011000101000",
2568 => "011011010110100000111010",
2569 => "011000110110101100111101",
2570 => "100010100111011101000101",
2571 => "010001010011000100011010",
2572 => "000101000000110000001011",
2573 => "000000000000000000000000",
2574 => "000000000000000000000000",
2575 => "000000000000000000000000",
2576 => "000000100000001000000010",
2577 => "001001110011010000101100",
2578 => "000110010010001000011100",
2579 => "000000000000000000000000",
2580 => "000000000000000000000000",
2581 => "000000000000000000000000",
2582 => "000000000000000000000000",
2583 => "000000000000000000000000",
2584 => "000000000000000000000000",
2585 => "000000000000000000000000",
2586 => "000000000000000000000000",
2587 => "000000000000000000000000",
2588 => "000000000000000000000000",
2589 => "000000000000000000000000",
2590 => "000000000000000000000000",
2591 => "000000000000000000000000",
2592 => "000000000000000000000000",
2593 => "000000000000000000000000",
2594 => "000000000000000000000000",
2595 => "000000000000000000000000",
2596 => "000000000000000000000000",
2597 => "000000000000000000000000",
2598 => "000000000000000000000000",
2599 => "000000000000000000000000",
2600 => "000000000000000000000000",
2601 => "000000000000000000000000",
2602 => "000000000000000000000000",
2603 => "000000000000000000000000",
2604 => "000000000000000000000000",
2605 => "000000000000000000000000",
2606 => "000000000000000000000000",
2607 => "000011100001001000001111",
2608 => "001101010100001000111100",
2609 => "000001000000010000000100",
2610 => "000000000000000000000000",
2611 => "000000000000000000000000",
2612 => "000000000000000000000000",
2613 => "001000010000111100001001",
2614 => "011001110010101100100000",
2615 => "011010000101100100110011",
2616 => "010010000100110000110010",
2617 => "011001000110000000111100",
2618 => "011001010010011000100001",
2619 => "001000010000111100001111",
2620 => "000001110000010000111110",
2621 => "000001100000001101101010",
2622 => "000001110000011101101101",
2623 => "010000000100100110101110",
2624 => "001101100100101110101110",
2625 => "001100100011101001111011",
2626 => "000011000000110100110100",
2627 => "000010110000110000011000",
2628 => "000011000001001100011000",
2629 => "000010110000101100101110",
2630 => "001100000011101001111110",
2631 => "001101100100100010101110",
2632 => "001111110100101110110001",
2633 => "000010010000011101101110",
2634 => "000001010000010001101101",
2635 => "000010010000010000111111",
2636 => "000111100000101100010010",
2637 => "011010110010011000011101",
2638 => "011001000101110000111110",
2639 => "010010010100110000110111",
2640 => "011001100101100100110101",
2641 => "011001010010100100011101",
2642 => "001000000000110000001011",
2643 => "000000000000000000000000",
2644 => "000000000000000000000000",
2645 => "000000000000000000000000",
2646 => "000001000000001100000011",
2647 => "001101010100000000111001",
2648 => "000011110001001000010000",
2649 => "000000000000000000000000",
2650 => "000000000000000000000000",
2651 => "000000000000000000000000",
2652 => "000000000000000000000000",
2653 => "000000000000000000000000",
2654 => "000000000000000000000000",
2655 => "000000000000000000000000",
2656 => "000000000000000000000000",
2657 => "000000000000000000000000",
2658 => "000000000000000000000000",
2659 => "000000000000000000000000",
2660 => "000000000000000000000000",
2661 => "000000000000000000000000",
2662 => "000000000000000000000000",
2663 => "000000000000000000000000",
2664 => "000000000000000000000000",
2665 => "000000000000000000000000",
2666 => "000000000000000000000000",
2667 => "000000000000000000000000",
2668 => "000000000000000000000000",
2669 => "000000000000000000000000",
2670 => "000000000000000000000000",
2671 => "000000000000000000000000",
2672 => "000000000000000000000000",
2673 => "000000000000000000000000",
2674 => "000000000000000000000000",
2675 => "000000000000000000000000",
2676 => "000000000000000000000000",
2677 => "000011100000111000001101",
2678 => "001011010011011100110000",
2679 => "000001010000010100000101",
2680 => "000000000000000000000000",
2681 => "000000000000000000000000",
2682 => "000000000000000000000000",
2683 => "000011010000101000000111",
2684 => "001011010010011000011001",
2685 => "011000010101100100111010",
2686 => "010101100101011000110101",
2687 => "100010100111101101000110",
2688 => "001100100010011000011001",
2689 => "000010010000100100011000",
2690 => "000001000000001100101010",
2691 => "000001100000001100111011",
2692 => "000001110000010101000110",
2693 => "000000110000010000100000",
2694 => "000001010000001100110111",
2695 => "000001000000011101011100",
2696 => "000001000000010101100001",
2697 => "000101110001111000101110",
2698 => "001001010011000101000110",
2699 => "000001100000010101001001",
2700 => "000001100000010001001000",
2701 => "000001000000010000101101",
2702 => "000001110000001100100000",
2703 => "000001000000010001001000",
2704 => "000001100000001100111010",
2705 => "000001100000001100100101",
2706 => "000010000000011100010111",
2707 => "001011010010010000011001",
2708 => "100010010111101001001010",
2709 => "010110110101100100110101",
2710 => "011000100101100100111000",
2711 => "001100010010011000010111",
2712 => "000011010000100100000110",
2713 => "000000000000000000000000",
2714 => "000000000000000000000000",
2715 => "000000000000000000000000",
2716 => "000001010000010000000100",
2717 => "001011000011011100101111",
2718 => "000011000000111000001101",
2719 => "000000000000000000000000",
2720 => "000000000000000000000000",
2721 => "000000000000000000000000",
2722 => "000000000000000000000000",
2723 => "000000000000000000000000",
2724 => "000000000000000000000000",
2725 => "000000000000000000000000",
2726 => "000000000000000000000000",
2727 => "000000000000000000000000",
2728 => "000000000000000000000000",
2729 => "000000000000000000000000",
2730 => "000000000000000000000000",
2731 => "000000000000000000000000",
2732 => "000000000000000000000000",
2733 => "000000000000000000000000",
2734 => "000000000000000000000000",
2735 => "000000000000000000000000",
2736 => "000000000000000000000000",
2737 => "000000000000000000000000",
2738 => "000000000000000000000000",
2739 => "000000000000000000000000",
2740 => "000000000000000000000000",
2741 => "000000000000000000000000",
2742 => "000000000000000000000000",
2743 => "000000000000000000000000",
2744 => "000000000000000000000000",
2745 => "000000000000000000000000",
2746 => "000000000000000000000000",
2747 => "000001110000100000000111",
2748 => "001001100011010000101100",
2749 => "000011110001001000010001",
2750 => "000000000000000000000000",
2751 => "000000000000000000000000",
2752 => "000000000000000000000000",
2753 => "000111010000111000001100",
2754 => "010101110010111100011110",
2755 => "100000110111001100111110",
2756 => "010110000101001000110011",
2757 => "011001100101110100110110",
2758 => "010100100010011000100010",
2759 => "000110110000110000100110",
2760 => "000001110000010101010011",
2761 => "000010000000001101111011",
2762 => "000001000000010001011001",
2763 => "000001010000010100111110",
2764 => "000010110000110000111000",
2765 => "000010110000101101011000",
2766 => "000011010000111001101101",
2767 => "001010000011010101000011",
2768 => "001101010100011101001110",
2769 => "000001100000011101000111",
2770 => "000011000000101101011000",
2771 => "000010010000110101011011",
2772 => "000000110000100100111100",
2773 => "000001010000001101011010",
2774 => "000001000000010001110101",
2775 => "000001010000010101010101",
2776 => "000101100000110000011111",
2777 => "010100110010010000100011",
2778 => "011010100101101000110101",
2779 => "010110110101011000111000",
2780 => "100000100111000101000010",
2781 => "010101110011000000011101",
2782 => "000111000000110100001100",
2783 => "000000000000000000000000",
2784 => "000000000000000000000000",
2785 => "000000000000000000000000",
2786 => "000010110000110100001011",
2787 => "001001100011010000101011",
2788 => "000001100000100000000110",
2789 => "000000000000000000000000",
2790 => "000000000000000000000000",
2791 => "000000000000000000000000",
2792 => "000000000000000000000000",
2793 => "000000000000000000000000",
2794 => "000000000000000000000000",
2795 => "000000000000000000000000",
2796 => "000000000000000000000000",
2797 => "000000000000000000000000",
2798 => "000000000000000000000000",
2799 => "000000000000000000000000",
2800 => "000000000000000000000000",
2801 => "000000000000000000000000",
2802 => "000000000000000000000000",
2803 => "000000000000000000000000",
2804 => "000000000000000000000000",
2805 => "000000000000000000000000",
2806 => "000000000000000000000000",
2807 => "000000000000000000000000",
2808 => "000000000000000000000000",
2809 => "000000000000000000000000",
2810 => "000000000000000000000000",
2811 => "000000000000000000000000",
2812 => "000000000000000000000000",
2813 => "000000000000000000000000",
2814 => "000000000000000000000000",
2815 => "000000000000000000000000",
2816 => "000000000000000000000000",
2817 => "000010110000110000001011",
2818 => "001110000100100001000000",
2819 => "000101000001101000010110",
2820 => "000000000000000000000000",
2821 => "000000000000000000000000",
2822 => "000000000000000000000000",
2823 => "000111110000111000001100",
2824 => "010111010010110100011110",
2825 => "011011110110011001000100",
2826 => "010001000100000100101011",
2827 => "011001000101110000111000",
2828 => "010101100010100000011100",
2829 => "001000000000111000011001",
2830 => "000000110000000100110001",
2831 => "000000010000001000111111",
2832 => "000001000000010001011110",
2833 => "000100100001000001010000",
2834 => "000010100000101100101110",
2835 => "000100010001000101001101",
2836 => "000101100010000001000100",
2837 => "001101000100101001000011",
2838 => "010001010110000101010101",
2839 => "000101110001111101001010",
2840 => "000100000001000001000110",
2841 => "000010100000110000101100",
2842 => "000010100000011100110100",
2843 => "000001100000010101001111",
2844 => "000000100000000101000100",
2845 => "000000110000001100101011",
2846 => "000110110000110000011001",
2847 => "010110100010100100011110",
2848 => "010111110101110000111011",
2849 => "010001110100000100100110",
2850 => "011011010110010001000001",
2851 => "010111000010111100011111",
2852 => "000111000000110100001100",
2853 => "000000000000000000000000",
2854 => "000000000000000000000000",
2855 => "000000000000000000000000",
2856 => "000100000001010100010001",
2857 => "001110000100100000111110",
2858 => "000010010000101000001001",
2859 => "000000000000000000000000",
2860 => "000000000000000000000000",
2861 => "000000000000000000000000",
2862 => "000000000000000000000000",
2863 => "000000000000000000000000",
2864 => "000000000000000000000000",
2865 => "000000000000000000000000",
2866 => "000000000000000000000000",
2867 => "000000000000000000000000",
2868 => "000000000000000000000000",
2869 => "000000000000000000000000",
2870 => "000000000000000000000000",
2871 => "000000000000000000000000",
2872 => "000000000000000000000000",
2873 => "000000000000000000000000",
2874 => "000000000000000000000000",
2875 => "000000000000000000000000",
2876 => "000000000000000000000000",
2877 => "000000000000000000000000",
2878 => "000000000000000000000000",
2879 => "000000000000000000000000",
2880 => "000000000000000000000000",
2881 => "000000000000000000000000",
2882 => "000000000000000000000000",
2883 => "000000000000000000000000",
2884 => "000000000000000000000000",
2885 => "000000000000000000000000",
2886 => "000000000000000000000000",
2887 => "000001110000011100000111",
2888 => "001001110011000100101010",
2889 => "000111110010001100011110",
2890 => "000000000000000000000000",
2891 => "000000000000000000000000",
2892 => "000000000000000000000000",
2893 => "000100000000100100001011",
2894 => "001010000010001000010101",
2895 => "010110110101010000110011",
2896 => "010100110100110000110000",
2897 => "011111110111001001000000",
2898 => "001010000010010000011100",
2899 => "001010010010001100111010",
2900 => "001010100010010001010100",
2901 => "000001010000010101001100",
2902 => "000001110000010101100100",
2903 => "000101010001011100110110",
2904 => "000110100001110001000111",
2905 => "000101100001101100111101",
2906 => "001010010011110001000010",
2907 => "001010000011110101000001",
2908 => "001100100100100001001101",
2909 => "001010110100110101010000",
2910 => "000111100010010001000110",
2911 => "000110100001101001000110",
2912 => "000101010001010100110100",
2913 => "000001010000011001100000",
2914 => "000001010000010001001111",
2915 => "001010010010011001010111",
2916 => "001010100010010100111111",
2917 => "001001010010001000010111",
2918 => "011111110110111001000101",
2919 => "010101000100111100101101",
2920 => "010110010101001100110110",
2921 => "001010000010010000010101",
2922 => "000011000000100000000110",
2923 => "000000000000000000000000",
2924 => "000000000000000000000000",
2925 => "000000000000000000000000",
2926 => "000110100001111000011001",
2927 => "001001000011001000101000",
2928 => "000001100000011100000110",
2929 => "000000000000000000000000",
2930 => "000000000000000000000000",
2931 => "000000000000000000000000",
2932 => "000000000000000000000000",
2933 => "000000000000000000000000",
2934 => "000000000000000000000000",
2935 => "000000000000000000000000",
2936 => "000000000000000000000000",
2937 => "000000000000000000000000",
2938 => "000000000000000000000000",
2939 => "000000000000000000000000",
2940 => "000000000000000000000000",
2941 => "000000000000000000000000",
2942 => "000000000000000000000000",
2943 => "000000000000000000000000",
2944 => "000000000000000000000000",
2945 => "000000000000000000000000",
2946 => "000000000000000000000000",
2947 => "000000000000000000000000",
2948 => "000000000000000000000000",
2949 => "000000000000000000000000",
2950 => "000000000000000000000000",
2951 => "000000000000000000000000",
2952 => "000000000000000000000000",
2953 => "000000000000000000000000",
2954 => "000000000000000000000000",
2955 => "000000000000000000000000",
2956 => "000000000000000000000000",
2957 => "000010010000101000001010",
2958 => "001110110100100101000001",
2959 => "001010000011000100101001",
2960 => "000000010000000100000001",
2961 => "000000000000000000000000",
2962 => "000000000000000000000000",
2963 => "001000010000110100001100",
2964 => "011000010011000100011111",
2965 => "100001110111011001000101",
2966 => "010111110101001000101101",
2967 => "011110100110101001000000",
2968 => "011000010101100100101110",
2969 => "011011010110000001000001",
2970 => "010110010101000000111111",
2971 => "000101000001001001000111",
2972 => "000010010000011001011011",
2973 => "001001010010111100101010",
2974 => "001100110100010100111111",
2975 => "001001110011010100101110",
2976 => "000110110011001001001000",
2977 => "000010110010010100110101",
2978 => "000001110001110000101111",
2979 => "000101110010111101000011",
2980 => "001011100100001000110110",
2981 => "001100100100011001000100",
2982 => "001001100011000100100111",
2983 => "000010000000011001011001",
2984 => "000101100001000001000110",
2985 => "010110000101000001000011",
2986 => "011010110110000001000000",
2987 => "011001000101100000110100",
2988 => "011110000110100000110110",
2989 => "010111110101100000110100",
2990 => "100001010111011001000001",
2991 => "011000110010111100011110",
2992 => "000111010000110000001010",
2993 => "000000000000000000000000",
2994 => "000000000000000000000000",
2995 => "000000000000000000000000",
2996 => "001000110010111100100110",
2997 => "001110100100101101000001",
2998 => "000010000000100100001000",
2999 => "000000000000000000000000",
3000 => "000000000000000000000000",
3001 => "000000000000000000000000",
3002 => "000000000000000000000000",
3003 => "000000000000000000000000",
3004 => "000000000000000000000000",
3005 => "000000000000000000000000",
3006 => "000000000000000000000000",
3007 => "000000000000000000000000",
3008 => "000000000000000000000000",
3009 => "000000000000000000000000",
3010 => "000000000000000000000000",
3011 => "000000000000000000000000",
3012 => "000000000000000000000000",
3013 => "000000000000000000000000",
3014 => "000000000000000000000000",
3015 => "000000000000000000000000",
3016 => "000000000000000000000000",
3017 => "000000000000000000000000",
3018 => "000000000000000000000000",
3019 => "000000000000000000000000",
3020 => "000000000000000000000000",
3021 => "000000000000000000000000",
3022 => "000000000000000000000000",
3023 => "000000000000000000000000",
3024 => "000000000000000000000000",
3025 => "000000000000000000000000",
3026 => "000000000000000000000000",
3027 => "000000010000000100000001",
3028 => "000110010010000000011010",
3029 => "001001000010111100100110",
3030 => "000010000000100000000111",
3031 => "000000000000000000000000",
3032 => "000000000000000000000000",
3033 => "000110010000101100001011",
3034 => "010011010010110100011011",
3035 => "011110110110110100111011",
3036 => "011010010101110000101111",
3037 => "011000010101011000110110",
3038 => "010101010100101100110010",
3039 => "010010000100000000101100",
3040 => "001100000010100100100100",
3041 => "000001100000011100100000",
3042 => "000001100000011001000110",
3043 => "000111010010011100100010",
3044 => "001010010011110100101111",
3045 => "001011100100001100111011",
3046 => "000111010011101101000101",
3047 => "000100100011010101010011",
3048 => "000100000011000000111101",
3049 => "000011010001010100010111",
3050 => "001100000100001100111011",
3051 => "001011000011110100101110",
3052 => "001000110010100000101000",
3053 => "000001000000010001000000",
3054 => "000001100000011000100100",
3055 => "001100000010011100100110",
3056 => "010011000011111000101001",
3057 => "010100110100100100110010",
3058 => "010111000101000100101101",
3059 => "011011010110000000111000",
3060 => "011110110110110000111010",
3061 => "010011010010110000100000",
3062 => "000101110000101000001001",
3063 => "000000000000000000000000",
3064 => "000000000000000000000000",
3065 => "000001100000010100000101",
3066 => "001001100010110100100101",
3067 => "000111010010000100011011",
3068 => "000000010000000100000001",
3069 => "000000000000000000000000",
3070 => "000000000000000000000000",
3071 => "000000000000000000000000",
3072 => "000000000000000000000000",
3073 => "000000000000000000000000",
3074 => "000000000000000000000000",
3075 => "000000000000000000000000",
3076 => "000000000000000000000000",
3077 => "000000000000000000000000",
3078 => "000000000000000000000000",
3079 => "000000000000000000000000",
3080 => "000000000000000000000000",
3081 => "000000000000000000000000",
3082 => "000000000000000000000000",
3083 => "000000000000000000000000",
3084 => "000000000000000000000000",
3085 => "000000000000000000000000",
3086 => "000000000000000000000000",
3087 => "000000000000000000000000",
3088 => "000000000000000000000000",
3089 => "000000000000000000000000",
3090 => "000000000000000000000000",
3091 => "000000000000000000000000",
3092 => "000000000000000000000000",
3093 => "000000000000000000000000",
3094 => "000000000000000000000000",
3095 => "000000000000000000000000",
3096 => "000000000000000000000000",
3097 => "000000010000000100000001",
3098 => "001001100010101100100111",
3099 => "001100010011111100110100",
3100 => "000101100001011100010101",
3101 => "000000000000000000000000",
3102 => "000000000000000000000000",
3103 => "000011000000100000000111",
3104 => "010010110100000000101010",
3105 => "011111000110110001000010",
3106 => "011000000101110100111100",
3107 => "001011000010111100100101",
3108 => "010011000100010000110000",
3109 => "010110110100111100111001",
3110 => "001011110010011100110000",
3111 => "000001110000011100111111",
3112 => "000001100000010101001101",
3113 => "000100010001010100011101",
3114 => "001010010011011000101000",
3115 => "001011000100001100111101",
3116 => "000100000010110000110100",
3117 => "000100000010011000110101",
3118 => "000101000011101001001001",
3119 => "000110100011101000111101",
3120 => "001011010100010000111001",
3121 => "001010010011011000101011",
3122 => "000101010001100000011101",
3123 => "000001000000010101000111",
3124 => "000001110000011001000000",
3125 => "001011110010010100101101",
3126 => "010110110100111000111011",
3127 => "010011110100011000110111",
3128 => "001001110011000000100001",
3129 => "011000000101101100111010",
3130 => "011110000110110101000010",
3131 => "010010100100001000101000",
3132 => "000010110000100000000101",
3133 => "000000000000000000000000",
3134 => "000000000000000000000000",
3135 => "000100010001001000010000",
3136 => "001100000011111000110100",
3137 => "001010000010111100101001",
3138 => "000000010000000100000001",
3139 => "000000000000000000000000",
3140 => "000000000000000000000000",
3141 => "000000000000000000000000",
3142 => "000000000000000000000000",
3143 => "000000000000000000000000",
3144 => "000000000000000000000000",
3145 => "000000000000000000000000",
3146 => "000000000000000000000000",
3147 => "000000000000000000000000",
3148 => "000000000000000000000000",
3149 => "000000000000000000000000",
3150 => "000000000000000000000000",
3151 => "000000000000000000000000",
3152 => "000000000000000000000000",
3153 => "000000000000000000000000",
3154 => "000000000000000000000000",
3155 => "000000000000000000000000",
3156 => "000000000000000000000000",
3157 => "000000000000000000000000",
3158 => "000000000000000000000000",
3159 => "000000000000000000000000",
3160 => "000000000000000000000000",
3161 => "000000000000000000000000",
3162 => "000000000000000000000000",
3163 => "000000000000000000000000",
3164 => "000000000000000000000000",
3165 => "000000000000000000000000",
3166 => "000000000000000000000000",
3167 => "000000000000000000000000",
3168 => "000101000001011100010100",
3169 => "001100110100000000110111",
3170 => "000101100001100100010100",
3171 => "000000000000000000000000",
3172 => "000000000000000000000000",
3173 => "000101110001010100010000",
3174 => "010101000101010000111001",
3175 => "010001110101000000111100",
3176 => "010000110110100101011011",
3177 => "001111010101000101001010",
3178 => "010100110100011100110100",
3179 => "010101110100110100111010",
3180 => "001100000010011000101110",
3181 => "000001010000010000110100",
3182 => "000001100000010001010010",
3183 => "000100110001010100011101",
3184 => "001011000011011100101111",
3185 => "001101000101011001001100",
3186 => "001011110110011101100000",
3187 => "000111100101111001010110",
3188 => "000111000101110001011100",
3189 => "001000100101010101010101",
3190 => "001100100101011101001010",
3191 => "001010110011100000110001",
3192 => "000101010001011100100010",
3193 => "000001110000001101010010",
3194 => "000001010000010000110011",
3195 => "001011100010010100101100",
3196 => "010110100100101100110110",
3197 => "010101100100100000110111",
3198 => "001110100100111101000100",
3199 => "010000100110101001011111",
3200 => "010001000101001100111001",
3201 => "010101000101001100111011",
3202 => "000101100001001100001110",
3203 => "000000000000000000000000",
3204 => "000000000000000000000000",
3205 => "000100110001010000010010",
3206 => "001100100011111100110110",
3207 => "000101010001101000010101",
3208 => "000000000000000000000000",
3209 => "000000000000000000000000",
3210 => "000000000000000000000000",
3211 => "000000000000000000000000",
3212 => "000000000000000000000000",
3213 => "000000000000000000000000",
3214 => "000000000000000000000000",
3215 => "000000000000000000000000",
3216 => "000000000000000000000000",
3217 => "000000000000000000000000",
3218 => "000000000000000000000000",
3219 => "000000000000000000000000",
3220 => "000000000000000000000000",
3221 => "000000000000000000000000",
3222 => "000000000000000000000000",
3223 => "000000000000000000000000",
3224 => "000000000000000000000000",
3225 => "000000000000000000000000",
3226 => "000000000000000000000000",
3227 => "000000000000000000000000",
3228 => "000000000000000000000000",
3229 => "000000000000000000000000",
3230 => "000000000000000000000000",
3231 => "000000000000000000000000",
3232 => "000000000000000000000000",
3233 => "000000000000000000000000",
3234 => "000000000000000000000000",
3235 => "000000000000000000000000",
3236 => "000000000000000000000000",
3237 => "000000010000000100000001",
3238 => "001000000010010100100000",
3239 => "001010010011100000101110",
3240 => "001011000011010100101110",
3241 => "000000010000000000000001",
3242 => "000000000000000000000000",
3243 => "000100010001001100010000",
3244 => "001110100101010101001000",
3245 => "010000010110100101100010",
3246 => "010000000110101001100010",
3247 => "001110010100011000111001",
3248 => "010000100011101000101011",
3249 => "011001100101001100111101",
3250 => "010000010011011100110100",
3251 => "000100010000110000101001",
3252 => "000001000000001100100100",
3253 => "000100100001010000010011",
3254 => "001001100011010100101011",
3255 => "001101100110011001010101",
3256 => "001010110110100101011011",
3257 => "001001010101100101010100",
3258 => "001000000101001101010110",
3259 => "001001110101011101010100",
3260 => "001110010110011101010011",
3261 => "001010010011010100101101",
3262 => "000101100001011100010101",
3263 => "000001000000001000100010",
3264 => "000100010000110000100100",
3265 => "010001010011010000110110",
3266 => "011000100101010000111001",
3267 => "010001000011110100101010",
3268 => "001111100011111100111000",
3269 => "010000010110100001100001",
3270 => "010000100110100101100001",
3271 => "001111010101001101001011",
3272 => "000100010001001000010000",
3273 => "000000000000000000000000",
3274 => "000000000000000000000000",
3275 => "001010010010111100101001",
3276 => "001010000011100000101101",
3277 => "001000010010100000100010",
3278 => "000000010000000100000001",
3279 => "000000000000000000000000",
3280 => "000000000000000000000000",
3281 => "000000000000000000000000",
3282 => "000000000000000000000000",
3283 => "000000000000000000000000",
3284 => "000000000000000000000000",
3285 => "000000000000000000000000",
3286 => "000000000000000000000000",
3287 => "000000000000000000000000",
3288 => "000000000000000000000000",
3289 => "000000000000000000000000",
3290 => "000000000000000000000000",
3291 => "000000000000000000000000",
3292 => "000000000000000000000000",
3293 => "000000000000000000000000",
3294 => "000000000000000000000000",
3295 => "000000000000000000000000",
3296 => "000000000000000000000000",
3297 => "000000000000000000000000",
3298 => "000000000000000000000000",
3299 => "000000000000000000000000",
3300 => "000000000000000000000000",
3301 => "000000000000000000000000",
3302 => "000000000000000000000000",
3303 => "000000000000000000000000",
3304 => "000000000000000000000000",
3305 => "000000000000000000000000",
3306 => "000000000000000000000000",
3307 => "000000010000000100000001",
3308 => "001000000010011100100000",
3309 => "001110110100101100111110",
3310 => "000111100010100000011110",
3311 => "000000100000001000000010",
3312 => "000000000000000000000000",
3313 => "000100000001001100010010",
3314 => "010000100110010101011100",
3315 => "010000000111000001101000",
3316 => "010000110101110001010111",
3317 => "011000010010000000100011",
3318 => "010011110010100000100010",
3319 => "011101100110011001000000",
3320 => "010100110100010000110110",
3321 => "001111000011000100101111",
3322 => "001000110001101100100100",
3323 => "000101010001001000010011",
3324 => "001000010010101100100011",
3325 => "001100100101010101001100",
3326 => "000111100100011001001000",
3327 => "000001100001001000100100",
3328 => "000010000001101100110001",
3329 => "000101010011110101000000",
3330 => "001011110101011001001001",
3331 => "001000110011000000100101",
3332 => "000100100000111100010011",
3333 => "001000010001101100100001",
3334 => "001110110011000000110010",
3335 => "010011110100010100110100",
3336 => "011101010110011101000001",
3337 => "010011100010011100011110",
3338 => "011000110010000000100111",
3339 => "010000000101100101001111",
3340 => "010000010110111001101001",
3341 => "001111100110011001011010",
3342 => "000011100001010000010001",
3343 => "000000000000000000000000",
3344 => "000000010000000100000000",
3345 => "000111100010001100011100",
3346 => "001110010100100000111011",
3347 => "001000110010101000100011",
3348 => "000000010000000100000001",
3349 => "000000000000000000000000",
3350 => "000000000000000000000000",
3351 => "000000000000000000000000",
3352 => "000000000000000000000000",
3353 => "000000000000000000000000",
3354 => "000000000000000000000000",
3355 => "000000000000000000000000",
3356 => "000000000000000000000000",
3357 => "000000000000000000000000",
3358 => "000000000000000000000000",
3359 => "000000000000000000000000",
3360 => "000000000000000000000000",
3361 => "000000000000000000000000",
3362 => "000000000000000000000000",
3363 => "000000000000000000000000",
3364 => "000000000000000000000000",
3365 => "000000000000000000000000",
3366 => "000000000000000000000000",
3367 => "000000000000000000000000",
3368 => "000000000000000000000000",
3369 => "000000000000000000000000",
3370 => "000000000000000000000000",
3371 => "000000000000000000000000",
3372 => "000000000000000000000000",
3373 => "000000000000000000000000",
3374 => "000000000000000000000000",
3375 => "000000000000000000000000",
3376 => "000000000000000000000000",
3377 => "000000000000000000000000",
3378 => "000101100001011100010010",
3379 => "001001110011000100100110",
3380 => "001001010010111000100011",
3381 => "000011000000110000001011",
3382 => "000000000000000000000000",
3383 => "000011100001001100010001",
3384 => "001111110110010001011011",
3385 => "010001000111001101101101",
3386 => "001111110110001001011101",
3387 => "010001010001110100011101",
3388 => "011011010011111100110100",
3389 => "011101110110100001000000",
3390 => "011001000101100000110111",
3391 => "010111010100111000110111",
3392 => "010100110100100100111010",
3393 => "001011100010011100100000",
3394 => "001001110011010000101101",
3395 => "001100000101011101001010",
3396 => "001010100110010001010110",
3397 => "000111100101011101010101",
3398 => "000110010100001101010011",
3399 => "001000110100111001010000",
3400 => "001100110101011001001001",
3401 => "001010000011011000110001",
3402 => "001010000010010000011101",
3403 => "010101000100101000110100",
3404 => "010111110100110100111010",
3405 => "011001100101011100110111",
3406 => "011101110110100100111101",
3407 => "011001000011110100110011",
3408 => "010010000001111000100000",
3409 => "001111100101111101010011",
3410 => "010001100111001001101100",
3411 => "001111100110010001011001",
3412 => "000011010001001000010000",
3413 => "000000000000000000000000",
3414 => "000010000000100000001000",
3415 => "001001100010111000100110",
3416 => "001001010011000100100111",
3417 => "000101110001100100010100",
3418 => "000000000000000000000000",
3419 => "000000000000000000000000",
3420 => "000000000000000000000000",
3421 => "000000000000000000000000",
3422 => "000000000000000000000000",
3423 => "000000000000000000000000",
3424 => "000000000000000000000000",
3425 => "000000000000000000000000",
3426 => "000000000000000000000000",
3427 => "000000000000000000000000",
3428 => "000000000000000000000000",
3429 => "000000000000000000000000",
3430 => "000000000000000000000000",
3431 => "000000000000000000000000",
3432 => "000000000000000000000000",
3433 => "000000000000000000000000",
3434 => "000000000000000000000000",
3435 => "000000000000000000000000",
3436 => "000000000000000000000000",
3437 => "000000000000000000000000",
3438 => "000000000000000000000000",
3439 => "000000000000000000000000",
3440 => "000000000000000000000000",
3441 => "000000000000000000000000",
3442 => "000000000000000000000000",
3443 => "000000000000000000000000",
3444 => "000000000000000000000000",
3445 => "000000000000000000000000",
3446 => "000000000000000000000000",
3447 => "000000000000000000000000",
3448 => "001000000010111000101001",
3449 => "001111100101100001001010",
3450 => "001001110011010100101010",
3451 => "000101100001011100010100",
3452 => "000000010000000100000001",
3453 => "000011000001000100010000",
3454 => "001111100110010001011010",
3455 => "010000110111001101101100",
3456 => "010001010111000001100110",
3457 => "001110110100100001000011",
3458 => "010011100100010100101011",
3459 => "011111000110101100111110",
3460 => "011100000110000000111001",
3461 => "011001100101001100111100",
3462 => "010110100100110000111010",
3463 => "001101000011000000100011",
3464 => "001010000011010100101111",
3465 => "001110110110000101010110",
3466 => "001010110110100001011000",
3467 => "001000100101001101010011",
3468 => "000100110011110001000011",
3469 => "001001010101001001001010",
3470 => "001110000110001001010001",
3471 => "001010010011100100110001",
3472 => "001100000010101100100000",
3473 => "010110100100110000110111",
3474 => "011001010101010000111001",
3475 => "011011100110000000111001",
3476 => "100000000110100000111011",
3477 => "010101110100101000101011",
3478 => "001111000100001100111110",
3479 => "010000010111000101100100",
3480 => "010001000111001101101100",
3481 => "001111100110001101011000",
3482 => "000011010001001000001111",
3483 => "000000000000000000000000",
3484 => "000100010001001100010000",
3485 => "001010100011011000101011",
3486 => "001111010101010101001000",
3487 => "001001100011001100101100",
3488 => "000000010000000100000001",
3489 => "000000000000000000000000",
3490 => "000000000000000000000000",
3491 => "000000000000000000000000",
3492 => "000000000000000000000000",
3493 => "000000000000000000000000",
3494 => "000000000000000000000000",
3495 => "000000000000000000000000",
3496 => "000000000000000000000000",
3497 => "000000000000000000000000",
3498 => "000000000000000000000000",
3499 => "000000000000000000000000",
3500 => "000000000000000000000000",
3501 => "000000000000000000000000",
3502 => "000000000000000000000000",
3503 => "000000000000000000000000",
3504 => "000000000000000000000000",
3505 => "000000000000000000000000",
3506 => "000000000000000000000000",
3507 => "000000000000000000000000",
3508 => "000000000000000000000000",
3509 => "000000000000000000000000",
3510 => "000000000000000000000000",
3511 => "000000000000000000000000",
3512 => "000000000000000000000000",
3513 => "000000000000000000000000",
3514 => "000000000000000000000000",
3515 => "000000000000000000000000",
3516 => "000000000000000000000000",
3517 => "000000000000000000000000",
3518 => "000011000000111100001110",
3519 => "001011100011110100110010",
3520 => "001001000010110100100010",
3521 => "000111100010000100011010",
3522 => "000011010000111000001100",
3523 => "000001110000100100001000",
3524 => "001110100101001001001100",
3525 => "001111110110101001100100",
3526 => "010000100110110001100011",
3527 => "010000110110101101100110",
3528 => "010011010101001100110111",
3529 => "100001000111001100111111",
3530 => "100011000111001101000001",
3531 => "011100110110010100111011",
3532 => "011001010101011000111001",
3533 => "010011110100010000110100",
3534 => "000111010010000000011100",
3535 => "001110110101110101010101",
3536 => "000111100100011001000101",
3537 => "000011010010110001001000",
3538 => "000011000010111101010000",
3539 => "000111000100000101000111",
3540 => "001111010101110001010010",
3541 => "000110100010010100011100",
3542 => "010011000100001100110100",
3543 => "011001000101010100110111",
3544 => "011101110110001100111001",
3545 => "100010110111001101000000",
3546 => "100000010111010001000010",
3547 => "010011100101011100110100",
3548 => "010001000110101001100011",
3549 => "001111110110110101100011",
3550 => "001111110110101001100100",
3551 => "001111000101010001001110",
3552 => "000010000000101000001001",
3553 => "000010000000100000000111",
3554 => "000110010001111100010111",
3555 => "001001100010110000100001",
3556 => "001011100011101100110000",
3557 => "000100000001010100010001",
3558 => "000000000000000000000000",
3559 => "000000000000000000000000",
3560 => "000000000000000000000000",
3561 => "000000000000000000000000",
3562 => "000000000000000000000000",
3563 => "000000000000000000000000",
3564 => "000000000000000000000000",
3565 => "000000000000000000000000",
3566 => "000000000000000000000000",
3567 => "000000000000000000000000",
3568 => "000000000000000000000000",
3569 => "000000000000000000000000",
3570 => "000000000000000000000000",
3571 => "000000000000000000000000",
3572 => "000000000000000000000000",
3573 => "000000000000000000000000",
3574 => "000000000000000000000000",
3575 => "000000000000000000000000",
3576 => "000000000000000000000000",
3577 => "000000000000000000000000",
3578 => "000000000000000000000000",
3579 => "000000000000000000000000",
3580 => "000000000000000000000000",
3581 => "000000000000000000000000",
3582 => "000000000000000000000000",
3583 => "000000000000000000000000",
3584 => "000000000000000000000000",
3585 => "000000000000000000000000",
3586 => "000000000000000000000000",
3587 => "000000000000000000000000",
3588 => "000101100001100100010101",
3589 => "001001000010111000100100",
3590 => "001010100011010100101001",
3591 => "001001100011001100100111",
3592 => "001001110011000100101010",
3593 => "000100000001000100010000",
3594 => "001001110011100100110101",
3595 => "010000100110111101100110",
3596 => "010000000110011101011111",
3597 => "010000100110111101100011",
3598 => "001111010101010001000111",
3599 => "010101100010111000100100",
3600 => "011100110010010000011100",
3601 => "011011110100110000110001",
3602 => "011101110110100000111101",
3603 => "011000110101011100111100",
3604 => "001000000010001000010111",
3605 => "001010000100111001000101",
3606 => "001001010110010001011111",
3607 => "000100010011101001001100",
3608 => "000011110010110101001000",
3609 => "001000010101101101011101",
3610 => "001010100101001001000110",
3611 => "000111100001111100010111",
3612 => "011000110101010100111011",
3613 => "011101110110011100111101",
3614 => "011011100100111000101111",
3615 => "011100010010010000100000",
3616 => "010101100010110100100011",
3617 => "001111010100111001000111",
3618 => "010000100110111001100101",
3619 => "010000000110100001011111",
3620 => "010000100110111101100110",
3621 => "001001110011100100110100",
3622 => "000011110000111100001111",
3623 => "001011100011000100101110",
3624 => "001001000011000000100110",
3625 => "001010100011010100100111",
3626 => "001001000010111100100010",
3627 => "000110110001101100010111",
3628 => "000000000000000000000000",
3629 => "000000000000000000000000",
3630 => "000000000000000000000000",
3631 => "000000000000000000000000",
3632 => "000000000000000000000000",
3633 => "000000000000000000000000",
3634 => "000000000000000000000000",
3635 => "000000000000000000000000",
3636 => "000000000000000000000000",
3637 => "000000000000000000000000",
3638 => "000000000000000000000000",
3639 => "000000000000000000000000",
3640 => "000000000000000000000000",
3641 => "000000000000000000000000",
3642 => "000000000000000000000000",
3643 => "000000000000000000000000",
3644 => "000000000000000000000000",
3645 => "000000000000000000000000",
3646 => "000000000000000000000000",
3647 => "000000000000000000000000",
3648 => "000000000000000000000000",
3649 => "000000000000000000000000",
3650 => "000000000000000000000000",
3651 => "000000000000000000000000",
3652 => "000000000000000000000000",
3653 => "000000000000000000000000",
3654 => "000000000000000000000000",
3655 => "000000000000000000000000",
3656 => "000000000000000000000000",
3657 => "000000000000000000000000",
3658 => "001000000010011000100011",
3659 => "001110110101000001000110",
3660 => "001011110100000000110110",
3661 => "001010010011010100101100",
3662 => "000111100010101100100100",
3663 => "000110110010001000100000",
3664 => "000011100001001100010010",
3665 => "010000100110011101011110",
3666 => "010000010110110001100101",
3667 => "010001100111001001101010",
3668 => "010000000100001001000010",
3669 => "010111010001001000011110",
3670 => "011101110001000000011111",
3671 => "010001110001001000011011",
3672 => "011111110111000001000011",
3673 => "011011010110000000111010",
3674 => "010011010100010000110010",
3675 => "001001010100001100111001",
3676 => "001011000110100101011111",
3677 => "000111110101011101011001",
3678 => "000100010011011001000110",
3679 => "001000010101101001011011",
3680 => "001000100100100100111100",
3681 => "010001110100001000101110",
3682 => "011100000101111000111100",
3683 => "011111100110111101000101",
3684 => "010001100001010000010111",
3685 => "011101000001000100100001",
3686 => "011000000001000100011111",
3687 => "010000000011101100111101",
3688 => "010000100111001101101001",
3689 => "010000000110110101100101",
3690 => "010000000110011101011111",
3691 => "000011000001000100010000",
3692 => "000110100010000000011110",
3693 => "000111110010101000100100",
3694 => "001010010011010100101101",
3695 => "001011110011111100110100",
3696 => "001110010101000001000100",
3697 => "001000100010100100100110",
3698 => "000000000000000000000000",
3699 => "000000000000000000000000",
3700 => "000000000000000000000000",
3701 => "000000000000000000000000",
3702 => "000000000000000000000000",
3703 => "000000000000000000000000",
3704 => "000000000000000000000000",
3705 => "000000000000000000000000",
3706 => "000000000000000000000000",
3707 => "000000000000000000000000",
3708 => "000000000000000000000000",
3709 => "000000000000000000000000",
3710 => "000000000000000000000000",
3711 => "000000000000000000000000",
3712 => "000000000000000000000000",
3713 => "000000000000000000000000",
3714 => "000000000000000000000000",
3715 => "000000000000000000000000",
3716 => "000000000000000000000000",
3717 => "000000000000000000000000",
3718 => "000000000000000000000000",
3719 => "000000000000000000000000",
3720 => "000000000000000000000000",
3721 => "000000000000000000000000",
3722 => "000000000000000000000000",
3723 => "000000000000000000000000",
3724 => "000000000000000000000000",
3725 => "000000000000000000000000",
3726 => "000000000000000100000000",
3727 => "000000000000000000000000",
3728 => "000001010000010100000101",
3729 => "001011000011011000101111",
3730 => "001011010011011000101110",
3731 => "000111110010011100100000",
3732 => "001000010011000000101001",
3733 => "001100110100001100111100",
3734 => "000010000000110000001001",
3735 => "001010100100000000111001",
3736 => "010001010111000001101000",
3737 => "010001010111010101101110",
3738 => "010000000011100100111011",
3739 => "010111110001000000011011",
3740 => "101000000010000100101010",
3741 => "010101110001100000011100",
3742 => "010100000100011100101010",
3743 => "011001100101100100111010",
3744 => "010011110100101000110110",
3745 => "001011100100111101000000",
3746 => "001001000100111001001010",
3747 => "000011110010011100110001",
3748 => "000010100010001001000010",
3749 => "001000010100110101010000",
3750 => "001101100101000101000010",
3751 => "010010110100011000110001",
3752 => "011001110101011000111100",
3753 => "010100000100011100101100",
3754 => "010110100001010100011001",
3755 => "101000100010001000101100",
3756 => "010111010001001000011110",
3757 => "001111100011010100111001",
3758 => "010010010111000101101100",
3759 => "010000100111000101101000",
3760 => "001010100100000100111100",
3761 => "000001110000100100001000",
3762 => "001100110100001100111100",
3763 => "001001000011000000101001",
3764 => "000111000010100000011111",
3765 => "001010100011011100101110",
3766 => "001010110011011100101110",
3767 => "000001110000100000000111",
3768 => "000000000000000000000000",
3769 => "000000000000000000000000",
3770 => "000000000000000000000000",
3771 => "000000000000000000000000",
3772 => "000000000000000000000000",
3773 => "000000000000000000000000",
3774 => "000000000000000000000000",
3775 => "000000000000000000000000",
3776 => "000000000000000000000000",
3777 => "000000000000000000000000",
3778 => "000000000000000000000000",
3779 => "000000000000000000000000",
3780 => "000000000000000000000000",
3781 => "000000000000000000000000",
3782 => "000000000000000000000000",
3783 => "000000000000000000000000",
3784 => "000000000000000000000000",
3785 => "000000000000000000000000",
3786 => "000000000000000000000000",
3787 => "000000000000000000000000",
3788 => "000000000000000000000000",
3789 => "000000000000000000000000",
3790 => "000000000000000000000000",
3791 => "000000000000000000000000",
3792 => "000000000000000000000000",
3793 => "000000000000000000000000",
3794 => "000000000000000000000000",
3795 => "000100100001010000010100",
3796 => "001101100100010001000000",
3797 => "001011000011110000110111",
3798 => "001000100010110000100111",
3799 => "000100010001100100010001",
3800 => "000110010010011000011101",
3801 => "001100000100000000111000",
3802 => "001000100011000000101001",
3803 => "001011010011110100110110",
3804 => "000101110001111000011011",
3805 => "000011000001000000001111",
3806 => "001111110110001101011011",
3807 => "010001010111001101101010",
3808 => "010000000110001001011000",
3809 => "001011100001111100011110",
3810 => "010001000001001000011001",
3811 => "001101110010111100101111",
3812 => "001101100100010101000001",
3813 => "001010000011010100101100",
3814 => "001001010010110000100011",
3815 => "001010000100100100111110",
3816 => "001010010110000001011011",
3817 => "000111010100010101000111",
3818 => "000011100010111101000010",
3819 => "001010000101111001011011",
3820 => "001010100100110000111111",
3821 => "001001000010110100100011",
3822 => "001001110011010100101000",
3823 => "001100010100100000111101",
3824 => "001101000011010000101110",
3825 => "010001110001000100011001",
3826 => "001011100001101100011100",
3827 => "001111110110000001010110",
3828 => "010000110111001001101000",
3829 => "001111110110011001011101",
3830 => "000011100001001100010010",
3831 => "000101010001110000011001",
3832 => "001011100011111000110110",
3833 => "001000100010110000100110",
3834 => "001100100100010000111011",
3835 => "000110100010011000011110",
3836 => "000100100001100000010010",
3837 => "001000010010101100100101",
3838 => "001011010011100000110110",
3839 => "001110000100001100111111",
3840 => "000100110001010000010100",
3841 => "000000000000000000000000",
3842 => "000000000000000000000000",
3843 => "000000000000000000000000",
3844 => "000000000000000000000000",
3845 => "000000000000000000000000",
3846 => "000000000000000000000000",
3847 => "000000000000000000000000",
3848 => "000000000000000000000000",
3849 => "000000000000000000000000",
3850 => "000000000000000000000000",
3851 => "000000000000000000000000",
3852 => "000000000000000000000000",
3853 => "000000000000000000000000",
3854 => "000000000000000000000000",
3855 => "000000000000000000000000",
3856 => "000000000000000000000000",
3857 => "000000000000000000000000",
3858 => "000000000000000000000000",
3859 => "000000000000000000000000",
3860 => "000000000000000000000000",
3861 => "000000000000000000000000",
3862 => "000000000000000000000000",
3863 => "000000000000000000000000",
3864 => "000000000000000000000000",
3865 => "000000000000000000000000",
3866 => "000000010000000100000001",
3867 => "000010110000111100001110",
3868 => "001110000100001100111110",
3869 => "001000010010101000100010",
3870 => "010001010101001101001010",
3871 => "001101010100011100111111",
3872 => "001000010011001000101001",
3873 => "001101000100101001000000",
3874 => "000110110010100100100100",
3875 => "000000000000000000000000",
3876 => "000100100001110000011010",
3877 => "010010110110111001100101",
3878 => "010001000110111101100011",
3879 => "010000000110011101011101",
3880 => "010000000110000101011000",
3881 => "001111110110011101011001",
3882 => "001110000101111001010111",
3883 => "001110100101111101010110",
3884 => "001110110101111001010100",
3885 => "001010000011101000110101",
3886 => "000011110001101100011010",
3887 => "001010110011101100111000",
3888 => "001011000011101000111001",
3889 => "000011110001011100010110",
3890 => "001001000011100000110000",
3891 => "001110100101111001010101",
3892 => "001110000110000001010110",
3893 => "001110100101111001010110",
3894 => "001111100110100001011010",
3895 => "010000110101111101011001",
3896 => "010000100110010101011010",
3897 => "010001010110111001100110",
3898 => "010011010110111101101000",
3899 => "000101100010000100011111",
3900 => "000000000000000000000000",
3901 => "000110110010011000100011",
3902 => "001101010100100100111111",
3903 => "001000010011001000100111",
3904 => "001100000100010000111011",
3905 => "010010110101010001001100",
3906 => "001000010010101000100010",
3907 => "001101000100001100111100",
3908 => "000011000001000100010000",
3909 => "000000010000000100000001",
3910 => "000000000000000000000000",
3911 => "000000000000000000000000",
3912 => "000000000000000000000000",
3913 => "000000000000000000000000",
3914 => "000000000000000000000000",
3915 => "000000000000000000000000",
3916 => "000000000000000000000000",
3917 => "000000000000000000000000",
3918 => "000000000000000000000000",
3919 => "000000000000000000000000",
3920 => "000000000000000000000000",
3921 => "000000000000000000000000",
3922 => "000000000000000000000000",
3923 => "000000000000000000000000",
3924 => "000000000000000000000000",
3925 => "000000000000000000000000",
3926 => "000000000000000000000000",
3927 => "000000000000000000000000",
3928 => "000000000000000000000000",
3929 => "000000000000000000000000",
3930 => "000000000000000000000000",
3931 => "000000000000000000000000",
3932 => "000000000000000000000000",
3933 => "000000000000000000000000",
3934 => "000000000000000000000000",
3935 => "000000000000000000000000",
3936 => "000001010000010100000101",
3937 => "000000100000001000000010",
3938 => "000101000001011100010100",
3939 => "001011000011101000110001",
3940 => "001000110010111100101000",
3941 => "010000100101000001001000",
3942 => "001100110100010100111011",
3943 => "001011100100001100111000",
3944 => "010000000101101101010010",
3945 => "000001010000011100000111",
3946 => "000000000000000000000000",
3947 => "000110000001110100011100",
3948 => "010100000110111101100101",
3949 => "010010100111011001101010",
3950 => "010011100111110001110010",
3951 => "010001000110101001100011",
3952 => "001110010101100101010011",
3953 => "001111010110000001011001",
3954 => "010010100111011001101100",
3955 => "010010100110111001100100",
3956 => "001011110100100001000000",
3957 => "001010110100000000111000",
3958 => "001011010011111000111001",
3959 => "001011100100010101000000",
3960 => "010010000110110001100011",
3961 => "010010110111100001101101",
3962 => "001111010110000101011010",
3963 => "001101100101100001010010",
3964 => "010000100110110001100011",
3965 => "010011010111101101110001",
3966 => "010010110111011001101010",
3967 => "010100000111000101100111",
3968 => "000110110010001100100001",
3969 => "000000000000000000000000",
3970 => "000001010000011100000111",
3971 => "001111010101100001010011",
3972 => "001011010100010100111000",
3973 => "001101000100010000110111",
3974 => "010000000101001001001011",
3975 => "001001010011000000101000",
3976 => "001010010011011100101110",
3977 => "000101110001100100010110",
3978 => "000000010000001000000010",
3979 => "000001010000010100000101",
3980 => "000000000000000000000000",
3981 => "000000000000000000000000",
3982 => "000000000000000000000000",
3983 => "000000000000000000000000",
3984 => "000000000000000000000000",
3985 => "000000000000000000000000",
3986 => "000000000000000000000000",
3987 => "000000000000000000000000",
3988 => "000000000000000000000000",
3989 => "000000000000000000000000",
3990 => "000000000000000000000000",
3991 => "000000000000000000000000",
3992 => "000000000000000000000000",
3993 => "000000000000000000000000",
3994 => "000000000000000000000000",
3995 => "000000000000000000000000",
3996 => "000000000000000000000000",
3997 => "000000000000000000000000",
3998 => "000000000000000000000000",
3999 => "000000000000000000000000",
4000 => "000000000000000000000000",
4001 => "000000000000000000000000",
4002 => "000000000000000000000000",
4003 => "000000000000000000000000",
4004 => "000000000000000000000000",
4005 => "000000000000000000000000",
4006 => "000110010001100100011010",
4007 => "001001000010110100101010",
4008 => "001100000100001000111010",
4009 => "001101100100110001000011",
4010 => "000101000010011000011110",
4011 => "001011100011110100110101",
4012 => "001010010011010000110000",
4013 => "001011010100010100111001",
4014 => "010001010110100101011011",
4015 => "000110000010000100011110",
4016 => "000000000000000000000000",
4017 => "000000000000000000000000",
4018 => "000101110010000000011100",
4019 => "010100100111001001100100",
4020 => "010110111000001101110111",
4021 => "010011000111010101101100",
4022 => "010000000110010001011101",
4023 => "001101100101010001001101",
4024 => "001101010101010001001010",
4025 => "001110100101100001001111",
4026 => "010001100110001001011010",
4027 => "001101110101000001001000",
4028 => "010000000101101101010001",
4029 => "010001010110001101011000",
4030 => "001111010101100001001111",
4031 => "001110000101010001001010",
4032 => "001101010101001101001101",
4033 => "001111100110001101011100",
4034 => "010010100111011001101100",
4035 => "010110111000001001110110",
4036 => "010101010111001101100110",
4037 => "000111100010011100100010",
4038 => "000000000000000000000000",
4039 => "000000000000000000000000",
4040 => "000110010010000100011111",
4041 => "010000110110101001011110",
4042 => "001011110100010100111011",
4043 => "001010000011001100101110",
4044 => "001010110100000100110111",
4045 => "000110000010010100100000",
4046 => "001100100100101001000000",
4047 => "001011110100010000111100",
4048 => "001000010010110000101010",
4049 => "000110000001100100011010",
4050 => "000000000000000000000000",
4051 => "000000000000000000000000",
4052 => "000000000000000000000000",
4053 => "000000000000000000000000",
4054 => "000000000000000000000000",
4055 => "000000000000000000000000",
4056 => "000000000000000000000000",
4057 => "000000000000000000000000",
4058 => "000000000000000000000000",
4059 => "000000000000000000000000",
4060 => "000000000000000000000000",
4061 => "000000000000000000000000",
4062 => "000000000000000000000000",
4063 => "000000000000000000000000",
4064 => "000000000000000000000000",
4065 => "000000000000000000000000",
4066 => "000000000000000000000000",
4067 => "000000000000000000000000",
4068 => "000000000000000000000000",
4069 => "000000000000000000000000",
4070 => "000000000000000000000000",
4071 => "000000000000000000000000",
4072 => "000000000000000000000000",
4073 => "000000000000000000000000",
4074 => "000000000000000000000000",
4075 => "000000000000000000000000",
4076 => "000000000000000000000000",
4077 => "000000010000000100000001",
4078 => "000101000001100100011000",
4079 => "001110110101100001010000",
4080 => "001111000101100101010000",
4081 => "001100100100101001000000",
4082 => "001111110101101101010010",
4083 => "001100110101000101000011",
4084 => "001011100100001100111000",
4085 => "000101010001110000011001",
4086 => "000000000000000000000000",
4087 => "000000000000000000000000",
4088 => "000100000001001000001111",
4089 => "001001110011011100101010",
4090 => "001101000100101000111011",
4091 => "010010110110110001100000",
4092 => "010010000110111001100110",
4093 => "001111010101110101010101",
4094 => "001110000101000101000111",
4095 => "001011010100011000111011",
4096 => "001100010100101000111110",
4097 => "001101000100110101000010",
4098 => "010001100110000001010101",
4099 => "001100010100110001000000",
4100 => "001100000100011000111011",
4101 => "001110000101000001000110",
4102 => "001110000101110101010101",
4103 => "010001110110111001100110",
4104 => "010011010110101101100001",
4105 => "001101000100101000111111",
4106 => "001001100011011100101011",
4107 => "000100110001011000010011",
4108 => "000000000000000000000000",
4109 => "000000000000000000000000",
4110 => "000101010001110000011001",
4111 => "001011110100001000111000",
4112 => "001100010100111001000011",
4113 => "001111010101101001010011",
4114 => "001101010100101001000000",
4115 => "001111000101100001010001",
4116 => "001111010101100101010000",
4117 => "000101000001101100011000",
4118 => "000000010000000100000001",
4119 => "000000000000000000000000",
4120 => "000000000000000000000000",
4121 => "000000000000000000000000",
4122 => "000000000000000000000000",
4123 => "000000000000000000000000",
4124 => "000000000000000000000000",
4125 => "000000000000000000000000",
4126 => "000000000000000000000000",
4127 => "000000000000000000000000",
4128 => "000000000000000000000000",
4129 => "000000000000000000000000",
4130 => "000000000000000000000000",
4131 => "000000000000000000000000",
4132 => "000000000000000000000000",
4133 => "000000000000000000000000",
4134 => "000000000000000000000000",
4135 => "000000000000000000000000",
4136 => "000000000000000000000000",
4137 => "000000000000000000000000",
4138 => "000000000000000000000000",
4139 => "000000000000000000000000",
4140 => "000000000000000000000000",
4141 => "000000000000000000000000",
4142 => "000000000000000000000000",
4143 => "000000000000000000000000",
4144 => "000000000000000000000000",
4145 => "000000000000000000000000",
4146 => "000000000000000000000000",
4147 => "000000000000000000000000",
4148 => "000011000000110100001101",
4149 => "001100100100101101000100",
4150 => "010100000111010101101101",
4151 => "001001110011101100110010",
4152 => "010011110111001001100110",
4153 => "001110010101100101001110",
4154 => "001001110011011000101100",
4155 => "000100000001010000010010",
4156 => "000000000000000000000000",
4157 => "000000000000000000000000",
4158 => "000110110001100100010110",
4159 => "001101010100001000111001",
4160 => "001100000100011100111010",
4161 => "001010110011111100110010",
4162 => "001001100011001100110000",
4163 => "001101110100110101000100",
4164 => "001110000101001001001101",
4165 => "001101100101010101001000",
4166 => "001111100110010001010111",
4167 => "001110010101011001001011",
4168 => "010010100110101001011111",
4169 => "001111110110010001011010",
4170 => "001101100101010101001000",
4171 => "001101110101010101001100",
4172 => "001100110100111001000101",
4173 => "001001100011001100101101",
4174 => "001011000011111000110000",
4175 => "001100100100010100111010",
4176 => "001101010100010100110111",
4177 => "000111000001110100011010",
4178 => "000000000000000000000000",
4179 => "000000000000000000000000",
4180 => "000100000001001100010001",
4181 => "001010010011011000101011",
4182 => "001110000101100001001101",
4183 => "010100000111010001101000",
4184 => "001001100011110000101110",
4185 => "010100100111001001101010",
4186 => "001101010100110101000111",
4187 => "000010110000110000001100",
4188 => "000000000000000000000000",
4189 => "000000000000000000000000",
4190 => "000000000000000000000000",
4191 => "000000000000000000000000",
4192 => "000000000000000000000000",
4193 => "000000000000000000000000",
4194 => "000000000000000000000000",
4195 => "000000000000000000000000",
4196 => "000000000000000000000000",
4197 => "000000000000000000000000",
4198 => "000000000000000000000000",
4199 => "000000000000000000000000",
4200 => "000000000000000000000000",
4201 => "000000000000000000000000",
4202 => "000000000000000000000000",
4203 => "000000000000000000000000",
4204 => "000000000000000000000000",
4205 => "000000000000000000000000",
4206 => "000000000000000000000000",
4207 => "000000000000000000000000",
4208 => "000000000000000000000000",
4209 => "000000000000000000000000",
4210 => "000000000000000000000000",
4211 => "000000000000000000000000",
4212 => "000000000000000000000000",
4213 => "000000000000000000000000",
4214 => "000000000000000000000000",
4215 => "000000000000000000000000",
4216 => "000000000000000000000000",
4217 => "000000000000000000000000",
4218 => "000000110000001100000011",
4219 => "000100100001011100010101",
4220 => "010000010110000101011000",
4221 => "010010010111000001100101",
4222 => "010011100111011001101110",
4223 => "001101010101001001000101",
4224 => "001001100010101100100111",
4225 => "000001000000010100000100",
4226 => "000000000000000000000000",
4227 => "000001000000001100000011",
4228 => "001100100010110000101100",
4229 => "001100000011010000110100",
4230 => "001101110100110101000011",
4231 => "001111010101011001001111",
4232 => "000100010001100100100111",
4233 => "001011010011011001110111",
4234 => "001101110100110101010010",
4235 => "001110010101010101001100",
4236 => "010011000110111101101011",
4237 => "010000110101111101010000",
4238 => "010101010111011001101010",
4239 => "010010110111000101101101",
4240 => "001110000101011101001100",
4241 => "001110000100110101010100",
4242 => "001100000011101001111011",
4243 => "000100000001100000101000",
4244 => "001111000101011001001011",
4245 => "001110000100111001000110",
4246 => "001011110011001000110101",
4247 => "001011110010110000101110",
4248 => "000000110000001100000011",
4249 => "000000000000000000000000",
4250 => "000001010000010100000101",
4251 => "001010000010110000100110",
4252 => "001101110101000001000101",
4253 => "010011010111011101101110",
4254 => "010001110110111101100100",
4255 => "010000100110010101011100",
4256 => "000100110001100100011000",
4257 => "000000110000001100000011",
4258 => "000000000000000000000000",
4259 => "000000000000000000000000",
4260 => "000000000000000000000000",
4261 => "000000000000000000000000",
4262 => "000000000000000000000000",
4263 => "000000000000000000000000",
4264 => "000000000000000000000000",
4265 => "000000000000000000000000",
4266 => "000000000000000000000000",
4267 => "000000000000000000000000",
4268 => "000000000000000000000000",
4269 => "000000000000000000000000",
4270 => "000000000000000000000000",
4271 => "000000000000000000000000",
4272 => "000000000000000000000000",
4273 => "000000000000000000000000",
4274 => "000000000000000000000000",
4275 => "000000000000000000000000",
4276 => "000000000000000000000000",
4277 => "000000000000000000000000",
4278 => "000000000000000000000000",
4279 => "000000000000000000000000",
4280 => "000000000000000000000000",
4281 => "000000000000000000000000",
4282 => "000000000000000000000000",
4283 => "000000000000000000000000",
4284 => "000000000000000000000000",
4285 => "000000000000000000000000",
4286 => "000000000000000000000000",
4287 => "000000000000000000000000",
4288 => "000000000000000000000000",
4289 => "000000000000000000000000",
4290 => "000110000010001100011111",
4291 => "010001000110000001010111",
4292 => "010000100101010001001000",
4293 => "001010000011001100100111",
4294 => "000011100000110100001111",
4295 => "000101100001100000011000",
4296 => "000110110010010100011101",
4297 => "001011000011100000101110",
4298 => "000101000001011100011010",
4299 => "000111100001110000101010",
4300 => "001011010011010000111001",
4301 => "001110010101010101001111",
4302 => "000010010000111001010000",
4303 => "001011100011011011011001",
4304 => "010101000110001011000000",
4305 => "001110010101010101011000",
4306 => "010110101000001001110011",
4307 => "010001000110000101010110",
4308 => "010111100111111001110010",
4309 => "010111111000010101111000",
4310 => "001110000101010001010110",
4311 => "010011110110010110110101",
4312 => "001101000011100111011111",
4313 => "000010010000111001010011",
4314 => "001110010101010001001111",
4315 => "001011000011011100111001",
4316 => "001000010001100100101000",
4317 => "000101010001011000011010",
4318 => "001010110011011000101011",
4319 => "000111000010010000011111",
4320 => "000101010001011100010111",
4321 => "000011110000111100010001",
4322 => "001001010011000100100111",
4323 => "001111100101010001000101",
4324 => "010010010101111001010101",
4325 => "000110110010010100100000",
4326 => "000000000000000000000000",
4327 => "000000000000000000000000",
4328 => "000000000000000000000000",
4329 => "000000000000000000000000",
4330 => "000000000000000000000000",
4331 => "000000000000000000000000",
4332 => "000000000000000000000000",
4333 => "000000000000000000000000",
4334 => "000000000000000000000000",
4335 => "000000000000000000000000",
4336 => "000000000000000000000000",
4337 => "000000000000000000000000",
4338 => "000000000000000000000000",
4339 => "000000000000000000000000",
4340 => "000000000000000000000000",
4341 => "000000000000000000000000",
4342 => "000000000000000000000000",
4343 => "000000000000000000000000",
4344 => "000000000000000000000000",
4345 => "000000000000000000000000",
4346 => "000000000000000000000000",
4347 => "000000000000000000000000",
4348 => "000000000000000000000000",
4349 => "000000000000000000000000",
4350 => "000000000000000000000000",
4351 => "000000000000000000000000",
4352 => "000000000000000000000000",
4353 => "000000000000000000000000",
4354 => "000000000000000000000000",
4355 => "000000000000000000000000",
4356 => "000000000000000000000000",
4357 => "000000000000000000000000",
4358 => "000000000000000000000000",
4359 => "000000000000000000000000",
4360 => "000001000000001100000010",
4361 => "001111100011101100101110",
4362 => "011011010101111100111110",
4363 => "011001010101010100110101",
4364 => "001101110011001100101010",
4365 => "001100110100000000111011",
4366 => "001101000100111101000010",
4367 => "001010010011101000101101",
4368 => "000110110010000000011010",
4369 => "001001110010001000100010",
4370 => "001101110011001100101111",
4371 => "001101100100110101000101",
4372 => "000110000010001100101011",
4373 => "001100010011011101111111",
4374 => "010010110100111011001100",
4375 => "001000000011000101011110",
4376 => "010101100111101001101110",
4377 => "010000000101101101010000",
4378 => "010111101000000001110010",
4379 => "010101110111110101110010",
4380 => "001000000011001001011011",
4381 => "010010100100100011001011",
4382 => "001110110100000010001010",
4383 => "000101100010000100101001",
4384 => "001110010100101001000011",
4385 => "001101100011001100110000",
4386 => "001011000010010000100101",
4387 => "000101010001111000010111",
4388 => "001010010011101100110001",
4389 => "001101000100110001000011",
4390 => "001101000100001000111010",
4391 => "001101100011010000101000",
4392 => "011000100101001100110101",
4393 => "011011100110000100111111",
4394 => "010000010011110100110000",
4395 => "000000100000001000000010",
4396 => "000000000000000000000000",
4397 => "000000000000000000000000",
4398 => "000000000000000000000000",
4399 => "000000000000000000000000",
4400 => "000000000000000000000000",
4401 => "000000000000000000000000",
4402 => "000000000000000000000000",
4403 => "000000000000000000000000",
4404 => "000000000000000000000000",
4405 => "000000000000000000000000",
4406 => "000000000000000000000000",
4407 => "000000000000000000000000",
4408 => "000000000000000000000000",
4409 => "000000000000000000000000",
4410 => "000000000000000000000000",
4411 => "000000000000000000000000",
4412 => "000000000000000000000000",
4413 => "000000000000000000000000",
4414 => "000000000000000000000000",
4415 => "000000000000000000000000",
4416 => "000000000000000000000000",
4417 => "000000000000000000000000",
4418 => "000000000000000000000000",
4419 => "000000000000000000000000",
4420 => "000000000000000000000000",
4421 => "000000000000000000000000",
4422 => "000000000000000000000000",
4423 => "000000000000000000000000",
4424 => "000000000000000000000000",
4425 => "000000000000000000000000",
4426 => "000000000000000000000000",
4427 => "000000000000000000000000",
4428 => "000000000000000000000000",
4429 => "000000000000000000000000",
4430 => "000100100001000100010010",
4431 => "000111100010000100011101",
4432 => "010010000100001000101100",
4433 => "010100000100110000110010",
4434 => "001100110100011000111010",
4435 => "010011110110111101100101",
4436 => "001110110101110001010100",
4437 => "001011100011111100110011",
4438 => "001010000011000000101000",
4439 => "001100000010101100100100",
4440 => "010010100011111000110100",
4441 => "001011100011110100110110",
4442 => "001101110101001001000111",
4443 => "000101010010000000100100",
4444 => "000011100001100000110101",
4445 => "001011110100010101000101",
4446 => "010010010110111101100101",
4447 => "001101000100111101000110",
4448 => "010010100110110101100001",
4449 => "010010100111000001100100",
4450 => "001100010100011101000110",
4451 => "000011110001101000110110",
4452 => "000100110001110100100100",
4453 => "001110000101000101000101",
4454 => "001011110011110000110100",
4455 => "010010010011110100110100",
4456 => "001101100010110000100110",
4457 => "001001000011000000100110",
4458 => "001011010011111000110101",
4459 => "001110000101101101001110",
4460 => "010011110110111101100111",
4461 => "001101000100011000111011",
4462 => "010011010100110000110011",
4463 => "010010000100010000101100",
4464 => "000111100010000100011011",
4465 => "000011100001000000001110",
4466 => "000000000000000000000000",
4467 => "000000000000000000000000",
4468 => "000000000000000000000000",
4469 => "000000000000000000000000",
4470 => "000000000000000000000000",
4471 => "000000000000000000000000",
4472 => "000000000000000000000000",
4473 => "000000000000000000000000",
4474 => "000000000000000000000000",
4475 => "000000000000000000000000",
4476 => "000000000000000000000000",
4477 => "000000000000000000000000",
4478 => "000000000000000000000000",
4479 => "000000000000000000000000",
4480 => "000000000000000000000000",
4481 => "000000000000000000000000",
4482 => "000000000000000000000000",
4483 => "000000000000000000000000",
4484 => "000000000000000000000000",
4485 => "000000000000000000000000",
4486 => "000000000000000000000000",
4487 => "000000000000000000000000",
4488 => "000000000000000000000000",
4489 => "000000000000000000000000",
4490 => "000000000000000000000000",
4491 => "000000000000000000000000",
4492 => "000000000000000000000000",
4493 => "000000000000000000000000",
4494 => "000000000000000000000000",
4495 => "000000000000000000000000",
4496 => "000000000000000000000000",
4497 => "000000000000000000000000",
4498 => "000000000000000000000000",
4499 => "000000000000000000000000",
4500 => "000010010000100100001001",
4501 => "000011100000111100010000",
4502 => "000110010001111000011100",
4503 => "001101000100110101000100",
4504 => "010001010110101101100001",
4505 => "010010000110011101011110",
4506 => "010101000111001001100101",
4507 => "001111000101011101001111",
4508 => "001001000011000100101010",
4509 => "010010000100000000101100",
4510 => "011010110101100100111101",
4511 => "010001000100001100110011",
4512 => "001011010011111100111011",
4513 => "001101010100110000111100",
4514 => "001111010101100001001111",
4515 => "001011100100001100111001",
4516 => "001101000100111001000110",
4517 => "001101000100100001000001",
4518 => "010000100101101101010011",
4519 => "001101010100111101000111",
4520 => "001011100100001000110101",
4521 => "001110110101100101010000",
4522 => "001101100100101101000100",
4523 => "001011100011111100110101",
4524 => "010001100100001100110110",
4525 => "011010110101101101000000",
4526 => "010011110100000100101111",
4527 => "001000110010111000100111",
4528 => "001110010101011001001111",
4529 => "010100110111001001100011",
4530 => "010010010110011101011100",
4531 => "010001010110101101100001",
4532 => "001101010100110101000100",
4533 => "000110010001110100011001",
4534 => "000011100001000000001111",
4535 => "000010000000100000001000",
4536 => "000000000000000000000000",
4537 => "000000000000000000000000",
4538 => "000000000000000000000000",
4539 => "000000000000000000000000",
4540 => "000000000000000000000000",
4541 => "000000000000000000000000",
4542 => "000000000000000000000000",
4543 => "000000000000000000000000",
4544 => "000000000000000000000000",
4545 => "000000000000000000000000",
4546 => "000000000000000000000000",
4547 => "000000000000000000000000",
4548 => "000000000000000000000000",
4549 => "000000000000000000000000",
4550 => "000000000000000000000000",
4551 => "000000000000000000000000",
4552 => "000000000000000000000000",
4553 => "000000000000000000000000",
4554 => "000000000000000000000000",
4555 => "000000000000000000000000",
4556 => "000000000000000000000000",
4557 => "000000000000000000000000",
4558 => "000000000000000000000000",
4559 => "000000000000000000000000",
4560 => "000000000000000000000000",
4561 => "000000000000000000000000",
4562 => "000000000000000000000000",
4563 => "000000000000000000000000",
4564 => "000000000000000000000000",
4565 => "000000000000000000000000",
4566 => "000000000000000000000000",
4567 => "000000000000000000000000",
4568 => "000000000000000000000000",
4569 => "000000000000000000000000",
4570 => "000000000000000000000000",
4571 => "000000000000000000000000",
4572 => "000000010000000100000001",
4573 => "000110100010000000011100",
4574 => "001100000100100100111100",
4575 => "001100110100111101000110",
4576 => "010100000111001101100100",
4577 => "010000000110001001011011",
4578 => "001011000011000000100010",
4579 => "011110110110110001000101",
4580 => "011011000101110000111100",
4581 => "000111100001100100010011",
4582 => "000100100001011000010100",
4583 => "001011100100000100110111",
4584 => "001101100101000001000100",
4585 => "000110100010001100100001",
4586 => "001000000010101100100010",
4587 => "001010110011100100110010",
4588 => "001100100100011000111011",
4589 => "000111110010101000100110",
4590 => "000110100010001000011110",
4591 => "001101110100111101000100",
4592 => "001011110100000000111000",
4593 => "000100100001101000010110",
4594 => "001000010001101000010101",
4595 => "011010000101110000111101",
4596 => "011111100110111001000110",
4597 => "001011100010111100100001",
4598 => "001111110101111101011001",
4599 => "010011110111001101100110",
4600 => "001101100100111001000101",
4601 => "001100100100100100111110",
4602 => "000110100010000100011110",
4603 => "000000010000000100000001",
4604 => "000000000000000000000000",
4605 => "000000000000000000000000",
4606 => "000000000000000000000000",
4607 => "000000000000000000000000",
4608 => "000000000000000000000000",
4609 => "000000000000000000000000",
4610 => "000000000000000000000000",
4611 => "000000000000000000000000",
4612 => "000000000000000000000000",
4613 => "000000000000000000000000",
4614 => "000000000000000000000000",
4615 => "000000000000000000000000",
4616 => "000000000000000000000000",
4617 => "000000000000000000000000",
4618 => "000000000000000000000000",
4619 => "000000000000000000000000",
4620 => "000000000000000000000000",
4621 => "000000000000000000000000",
4622 => "000000000000000000000000",
4623 => "000000000000000000000000",
4624 => "000000000000000000000000",
4625 => "000000000000000000000000",
4626 => "000000000000000000000000",
4627 => "000000000000000000000000",
4628 => "000000000000000000000000",
4629 => "000000000000000000000000",
4630 => "000000000000000000000000",
4631 => "000000000000000000000000",
4632 => "000000000000000000000000",
4633 => "000000000000000000000000",
4634 => "000000000000000000000000",
4635 => "000000000000000000000000",
4636 => "000000000000000000000000",
4637 => "000000000000000000000000",
4638 => "000000000000000000000000",
4639 => "000000000000000000000000",
4640 => "000000000000000000000000",
4641 => "000000000000000000000000",
4642 => "000000000000000000000000",
4643 => "000000110000001100000011",
4644 => "001000100010111000100110",
4645 => "001101110101001101001010",
4646 => "001110110101100101010000",
4647 => "000111010010100100100110",
4648 => "010101000100101100111010",
4649 => "010010010100000000101001",
4650 => "000101010001001000001011",
4651 => "000000010000000000000000",
4652 => "000110100001111100011011",
4653 => "001010110011010000101101",
4654 => "001011110011100100110001",
4655 => "000100010001001100001111",
4656 => "000111110010101000011111",
4657 => "001100000100001000111000",
4658 => "001011110100000100110111",
4659 => "001000010010100000100001",
4660 => "000011100001000100001100",
4661 => "001011010011101100110010",
4662 => "001010100011010000101100",
4663 => "000110010010001000011101",
4664 => "000000010000000100000001",
4665 => "000101010001001000001101",
4666 => "010001110011111000101000",
4667 => "010110010101000100111100",
4668 => "000111100010100000100101",
4669 => "001110010101100001001110",
4670 => "001101100101010101001010",
4671 => "001000000010101000100101",
4672 => "000000100000001000000010",
4673 => "000000000000000000000000",
4674 => "000000000000000000000000",
4675 => "000000000000000000000000",
4676 => "000000000000000000000000",
4677 => "000000000000000000000000",
4678 => "000000000000000000000000",
4679 => "000000000000000000000000",
4680 => "000000000000000000000000",
4681 => "000000000000000000000000",
4682 => "000000000000000000000000",
4683 => "000000000000000000000000",
4684 => "000000000000000000000000",
4685 => "000000000000000000000000",
4686 => "000000000000000000000000",
4687 => "000000000000000000000000",
4688 => "000000000000000000000000",
4689 => "000000000000000000000000",
4690 => "000000000000000000000000",
4691 => "000000000000000000000000",
4692 => "000000000000000000000000",
4693 => "000000000000000000000000",
4694 => "000000000000000000000000",
4695 => "000000000000000000000000",
4696 => "000000000000000000000000",
4697 => "000000000000000000000000",
4698 => "000000000000000000000000",
4699 => "000000000000000000000000",
4700 => "000000000000000000000000",
4701 => "000000000000000000000000",
4702 => "000000000000000000000000",
4703 => "000000000000000000000000",
4704 => "000000000000000000000000",
4705 => "000000000000000000000000",
4706 => "000000000000000000000000",
4707 => "000000000000000000000000",
4708 => "000000000000000000000000",
4709 => "000000000000000000000000",
4710 => "000000000000000000000000",
4711 => "000000000000000000000000",
4712 => "000000000000000000000000",
4713 => "000000000000000000000000",
4714 => "000001000000010000000100",
4715 => "000010110000110100001100",
4716 => "000011010001000000010000",
4717 => "000111000001100000011101",
4718 => "000100000000110000001011",
4719 => "000000010000000100000001",
4720 => "000000000000000000000000",
4721 => "000000010000001000000010",
4722 => "001011100011100000110100",
4723 => "000011000001000100001101",
4724 => "001000110010111000101000",
4725 => "000011110001011100010010",
4726 => "001001110011000100101010",
4727 => "000110000001110100011001",
4728 => "000101000001100100010111",
4729 => "001001010010100100100110",
4730 => "000100010001100000010011",
4731 => "001001010010111100101001",
4732 => "000010110001000000001101",
4733 => "001011010011011100110100",
4734 => "000000110000001100000011",
4735 => "000000000000000000000000",
4736 => "000000010000000100000001",
4737 => "000011100000110000001011",
4738 => "000110110001100000011101",
4739 => "000011010001000000001111",
4740 => "000010010000110000001010",
4741 => "000000100000001000000010",
4742 => "000000000000000000000000",
4743 => "000000000000000000000000",
4744 => "000000000000000000000000",
4745 => "000000000000000000000000",
4746 => "000000000000000000000000",
4747 => "000000000000000000000000",
4748 => "000000000000000000000000",
4749 => "000000000000000000000000",
4750 => "000000000000000000000000",
4751 => "000000000000000000000000",
4752 => "000000000000000000000000",
4753 => "000000000000000000000000",
4754 => "000000000000000000000000",
4755 => "000000000000000000000000",
4756 => "000000000000000000000000",
4757 => "000000000000000000000000",
4758 => "000000000000000000000000",
4759 => "000000000000000000000000",
4760 => "000000000000000000000000",
4761 => "000000000000000000000000",
4762 => "000000000000000000000000",
4763 => "000000000000000000000000",
4764 => "000000000000000000000000",
4765 => "000000000000000000000000",
4766 => "000000000000000000000000",
4767 => "000000000000000000000000",
4768 => "000000000000000000000000",
4769 => "000000000000000000000000",
4770 => "000000000000000000000000",
4771 => "000000000000000000000000",
4772 => "000000000000000000000000",
4773 => "000000000000000000000000",
4774 => "000000000000000000000000",
4775 => "000000000000000000000000",
4776 => "000000000000000000000000",
4777 => "000000000000000000000000",
4778 => "000000000000000000000000",
4779 => "000000000000000000000000",
4780 => "000000000000000000000000",
4781 => "000000000000000000000000",
4782 => "000000000000000000000000",
4783 => "000000000000000000000000",
4784 => "000000000000000000000000",
4785 => "000000000000000000000000",
4786 => "000000000000000000000000",
4787 => "000000000000000000000000",
4788 => "000000000000000000000000",
4789 => "000000000000000000000000",
4790 => "000000000000000000000000",
4791 => "000010100000101000001011",
4792 => "000111100010010100100101",
4793 => "000010100000100100001010",
4794 => "000111110001111100100001",
4795 => "000001000000010000000101",
4796 => "000001010000010100000101",
4797 => "000000000000000000000000",
4798 => "000000000000000000000000",
4799 => "000001000000001100000100",
4800 => "000000110000010000000100",
4801 => "000110000001101000011010",
4802 => "000001100000011000000111",
4803 => "000110110010000000100000",
4804 => "000011000000110000001101",
4805 => "000000000000000000000000",
4806 => "000000000000000000000000",
4807 => "000000000000000000000000",
4808 => "000000000000000000000000",
4809 => "000000000000000000000000",
4810 => "000000000000000000000000",
4811 => "000000000000000000000000",
4812 => "000000000000000000000000",
4813 => "000000000000000000000000",
4814 => "000000000000000000000000",
4815 => "000000000000000000000000",
4816 => "000000000000000000000000",
4817 => "000000000000000000000000",
4818 => "000000000000000000000000",
4819 => "000000000000000000000000",
4820 => "000000000000000000000000",
4821 => "000000000000000000000000",
4822 => "000000000000000000000000",
4823 => "000000000000000000000000",
4824 => "000000000000000000000000",
4825 => "000000000000000000000000",
4826 => "000000000000000000000000",
4827 => "000000000000000000000000",
4828 => "000000000000000000000000",
4829 => "000000000000000000000000",
4830 => "000000000000000000000000",
4831 => "000000000000000000000000",
4832 => "000000000000000000000000",
4833 => "000000000000000000000000",
4834 => "000000000000000000000000",
4835 => "000000000000000000000000",
4836 => "000000000000000000000000",
4837 => "000000000000000000000000",
4838 => "000000000000000000000000",
4839 => "000000000000000000000000",
4840 => "000000000000000000000000",
4841 => "000000000000000000000000",
4842 => "000000000000000000000000",
4843 => "000000000000000000000000",
4844 => "000000000000000000000000",
4845 => "000000000000000000000000",
4846 => "000000000000000000000000",
4847 => "000000000000000000000000",
4848 => "000000000000000000000000",
4849 => "000000000000000000000000",
4850 => "000000000000000000000000",
4851 => "000000000000000000000000",
4852 => "000000000000000000000000",
4853 => "000000000000000000000000",
4854 => "000000000000000000000000",
4855 => "000000000000000000000000",
4856 => "000000000000000000000000",
4857 => "000000000000000000000000",
4858 => "000000000000000000000000",
4859 => "000000000000000000000000",
4860 => "000000000000000000000000",
4861 => "000000100000001000000010",
4862 => "000000100000000100000010",
4863 => "000000000000000000000000",
4864 => "000000000000000000000000",
4865 => "000000000000000000000000",
4866 => "000000000000000000000000",
4867 => "000000000000000000000000",
4868 => "000000000000000000000000",
4869 => "000000000000000000000000",
4870 => "000000000000000000000000",
4871 => "000000000000000000000000",
4872 => "000000000000000000000000",
4873 => "000000010000000100000001",
4874 => "000000100000001000000010",
4875 => "000000000000000000000000",
4876 => "000000000000000000000000",
4877 => "000000000000000000000000",
4878 => "000000000000000000000000",
4879 => "000000000000000000000000",
4880 => "000000000000000000000000",
4881 => "000000000000000000000000",
4882 => "000000000000000000000000",
4883 => "000000000000000000000000",
4884 => "000000000000000000000000",
4885 => "000000000000000000000000",
4886 => "000000000000000000000000",
4887 => "000000000000000000000000",
4888 => "000000000000000000000000",
4889 => "000000000000000000000000",
4890 => "000000000000000000000000",
4891 => "000000000000000000000000",
4892 => "000000000000000000000000",
4893 => "000000000000000000000000",
4894 => "000000000000000000000000",
4895 => "000000000000000000000000",
4896 => "000000000000000000000000",
4897 => "000000000000000000000000",
4898 => "000000000000000000000000",
4899 => "000000000000000000000000"

    );
begin
    data_out <= ROM_Data(to_integer(unsigned(address)));
end architecture Behavioral;