// PLL.v

// Generated using ACDS version 13.1 162 at 2024.05.17.15:27:36

`timescale 1 ps / 1 ps
module PLL (
		input  wire  clk_in_clk,  //  clk_in.clk
		input  wire  reset_reset, //   reset.reset
		output wire  clk_out_clk  // clk_out.clk
	);

	PLL_pll_0 pll_0 (
		.refclk   (clk_in_clk),  //  refclk.clk
		.rst      (reset_reset), //   reset.reset
		.outclk_0 (clk_out_clk), // outclk0.clk
		.locked   ()             // (terminated)
	);

endmodule
